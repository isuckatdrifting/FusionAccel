`timescale 1ns/1ps
// `define CMAC
// `define SACC
`define SCMP

module engine_tb;

reg 		clk;
//Control signals csb->engine
reg 		rst;
reg 		engine_valid;
reg [2:0] 	op_type;
reg	[3:0]	stride;
reg [15:0]  stride2;
reg [7:0]  	kernel;
reg [7:0]	kernel_size;
reg [15:0]  i_channel;
reg [15:0]  o_channel;
reg [7:0]	i_side;
reg [7:0]   o_side;
reg	[15:0]  bias;
//Response signals engine->csb
wire		gemm_finish;
//Command path engine->dma
wire        output_en;
wire [9:0]  d_ram_read_addr;
wire [12:0] w_ram_read_addr;
//Data path dma->engine
reg [127:0] input_data;
reg [127:0] input_weig;
//Data path engine->dma
wire [15:0]	output_data;

`ifdef CMAC
	reg [15:0] data [0:2783];
	reg [15:0] weight [0:1151];
	initial begin
	/*
	data[0] = 16'h4d86; data[1] = 16'h4cbd; data[2] = 16'h4a18; data[3] = 16'h0000; data[4] = 16'h4b7c; data[5] = 16'h4269; data[6] = 16'h59b9; data[7] = 16'h4d2f; data[8] = 16'h480c; data[9] = 16'h449a; data[10] = 16'h4e77; data[11] = 16'h37b9; data[12] = 16'h530a; data[13] = 16'h4d34; data[14] = 16'h4873; data[15] =
16'h4cb6; data[16] = 16'h0000; data[17] = 16'h45ee; data[18] = 16'h4c48; data[19] = 16'h4bea; data[20] = 16'h4bd0; data[21] = 16'h0000; data[22] = 16'h0000; data[23] = 16'h4ae0; data[24] = 16'h4c07; data[25] = 16'h4df6; data[26] = 16'h52ae; data[27] = 16'h4262; data[28] = 16'h5403; data[29] = 16'h0000; data[30] = 16'h4a2d; data[31] = 16'h5170; data[32] = 16'h4d30; data[33] = 16'h0000; data[34] = 16'h4843; data[35] = 16'h0000; data[36] = 16'h4604; data[37] = 16'h2871; data[38] = 16'h0000; data[39] = 16'h0000; data[40] = 16'h4e4f; data[41] = 16'h4cb8; data[42] = 16'h4c8c; data[43] = 16'h504d; data[44] = 16'h4e9d; data[45] = 16'h3660; data[46] = 16'h0000; data[47] = 16'h4908; data[48] = 16'h4ef9; data[49] = 16'h53c6; data[50] = 16'h472a; data[51] = 16'h58e1; data[52] = 16'h4b5c; data[53] = 16'h4910; data[54] = 16'h5049; data[55] = 16'h5411; data[56] = 16'h0000; data[57] = 16'h4fdf; data[58] = 16'h48a0; data[59] = 16'h4a80; data[60] = 16'h4e60; data[61] = 16'h4ab3; data[62] = 16'h4caa; data[63] = 16'h514c;

weight[0] = 16'h27ae; weight[1] = 16'had60; weight[2] = 16'h2dbf; weight[3] = 16'ha8b9; weight[4] = 16'h36db; weight[5] = 16'h2a8e; weight[6] = 16'h278d; weight[7] = 16'h3131; weight[8] = 16'hb2d8; weight[9] = 16'h2694; weight[10] = 16'hb4f5; weight[11] = 16'h35fd; weight[12] = 16'h26bc; weight[13] = 16'h28d0; weight[14] = 16'h2d8c; weight[15] = 16'hb44e; weight[16] = 16'h341c; weight[17] = 16'haef2; weight[18] = 16'h3420; weight[19] = 16'hb381; weight[20] = 16'h36e5; weight[21] = 16'h289f; weight[22] = 16'h2c19; weight[23] = 16'hac9a; weight[24]
= 16'hb32f; weight[25] = 16'h37a3; weight[26] = 16'h2c55; weight[27] = 16'h360e; weight[28] = 16'ha8fe; weight[29] = 16'ha93f; weight[30] = 16'hacf6; weight[31] = 16'hb0a9; weight[32] = 16'hb61e; weight[33] = 16'h31a2; weight[34] = 16'hb10f; weight[35] = 16'h349e; weight[36] = 16'h31cf; weight[37] = 16'hb4e5; weight[38] = 16'h2b5f; weight[39] = 16'h1cb6; weight[40] = 16'hb75f; weight[41] = 16'hb497; weight[42] = 16'h3197; weight[43] = 16'hb5b3; weight[44] = 16'hb64d; weight[45] = 16'h3683; weight[46] = 16'hb630; weight[47] = 16'h2ebd; weight[48] = 16'h3867; weight[49] = 16'h3118; weight[50] = 16'h23c8; weight[51] = 16'h2e77; weight[52] = 16'haf54; weight[53] = 16'hb622; weight[54] = 16'hb3e9; weight[55] = 16'h3471; weight[56] = 16'haa2b; weight[57] = 16'h353f; weight[58] = 16'h2a81; weight[59] = 16'h352e; weight[60] = 16'h3049; weight[61] = 16'h38ed; weight[62] = 16'ha9c9; weight[63] = 16'hb64f;*/
	/*
	data[0] = 16'hce83; data[1] = 16'h4f98; data[2] = 16'h4e17; data[3] = 16'h0000; 
	data[4] = 16'h0000; data[5] = 16'h0000; data[6] = 16'h0000; data[7] = 16'h0000; 
	data[8] = 16'hce24; data[9] = 16'h5087; data[10] = 16'h4F8D; data[11] = 16'h0000; 
	data[12] = 16'h0000; data[13] = 16'h0000; data[14] = 16'h0000; data[15] = 16'h0000; 
	data[16] = 16'hCCEF; data[17] = 16'h51FB; data[18] = 16'h50DE; data[19] = 16'h0000;
	data[20] = 16'h0000; data[21] = 16'h0000; data[22] = 16'h0000; data[23] = 16'h0000;

	data[24] = 16'hCDE5; data[25] = 16'h5087; data[26] = 16'h4F10; data[27] = 16'h0000; 
	data[28] = 16'h0000; data[29] = 16'h0000; data[30] = 16'h0000; data[31] = 16'h0000; 
	data[32] = 16'hCFEB; data[33] = 16'h4FA7; data[34] = 16'h4DA9; data[35] = 16'h0000; 
	data[36] = 16'h0000; data[37] = 16'h0000; data[38] = 16'h0000; data[39] = 16'h0000;
	data[40] = 16'hD035; data[41] = 16'h5050; data[42] = 16'h4E61; data[43] = 16'h0000; 
	data[44] = 16'h0000; data[45] = 16'h0000; data[46] = 16'h0000; data[47] = 16'h0000;

	data[48] = 16'hD0A0; data[49] = 16'h4E32; data[50] = 16'h4C33; data[51] = 16'h0000; 
	data[52] = 16'h0000; data[53] = 16'h0000; data[54] = 16'h0000; data[55] = 16'h0000; 
	data[56] = 16'hD151; data[57] = 16'h4D6D; data[58] = 16'h49E7; data[59] = 16'h0000;
	data[60] = 16'h0000; data[61] = 16'h0000; data[62] = 16'h0000; data[63] = 16'h0000; 
	data[64] = 16'hD157; data[65] = 16'h4E9C; data[66] = 16'h4BC3; data[67] = 16'h0000; 
	data[68] = 16'h0000; data[69] = 16'h0000; data[70] = 16'h0000; data[71] = 16'h0000; 
	
	data[72] = 16'hd2b2; data[73] = 16'h4bef; data[74] = 16'h405e; data[75] = 16'h0000; 
	data[76] = 16'h0000; data[77] = 16'h0000; data[78] = 16'h0000; data[79] = 16'h0000; 
	data[80] = 16'hd1fc; data[81] = 16'h4d8b; data[82] = 16'h482d; data[83] = 16'h0000;
	data[84] = 16'h0000; data[85] = 16'h0000; data[86] = 16'h0000; data[87] = 16'h0000; 
	data[88] = 16'hd1db; data[89] = 16'h4e52; data[90] = 16'h49b4; data[91] = 16'h0000;
	data[92] = 16'h0000; data[93] = 16'h0000; data[94] = 16'h0000; data[95] = 16'h0000; 

	data[96] = 16'hd37e; data[97] = 16'h4bba; data[98] = 16'h387c; data[99] = 16'h0000;
	data[100] = 16'h0000; data[101] = 16'h0000; data[102] = 16'h0000; data[103] = 16'h0000; 
	data[104] = 16'hd34c; data[105] = 16'h4c67; data[106] = 16'h414e; data[107] = 16'h0000;
	data[108] = 16'h0000; data[109] = 16'h0000; data[110] = 16'h0000; data[111] = 16'h0000; 
	data[112] = 16'hd2d5; data[113] = 16'h4cad; data[114] = 16'h44ab; data[115] = 16'h0000;
	data[116] = 16'h0000; data[117] = 16'h0000; data[118] = 16'h0000; data[119] = 16'h0000; 

	data[120] = 16'hd43b; data[121] = 16'h480b; data[122] = 16'hc7ca; data[123] = 16'h0000;
	data[124] = 16'h0000; data[125] = 16'h0000; data[126] = 16'h0000; data[127] = 16'h0000; 
	data[128] = 16'hd453; data[129] = 16'h472b; data[130] = 16'hc863; data[131] = 16'h0000;
	data[132] = 16'h0000; data[133] = 16'h0000; data[134] = 16'h0000; data[135] = 16'h0000; 
	data[136] = 16'hd30c; data[137] = 16'h4c7e; data[138] = 16'h4030; data[139] = 16'h0000;
	data[140] = 16'h0000; data[141] = 16'h0000; data[142] = 16'h0000; data[143] = 16'h0000;

	data[144] = 16'hd29a; data[145] = 16'h4c60; data[146] = 16'h40ea; data[147] = 16'h0000;
	data[148] = 16'h0000; data[149] = 16'h0000; data[150] = 16'h0000; data[151] = 16'h0000;
	data[152] = 16'hd2ce; data[153] = 16'h4b51; data[154] = 16'hb765; data[155] = 16'h0000;
	data[156] = 16'h0000; data[157] = 16'h0000; data[158] = 16'h0000; data[159] = 16'h0000;
	data[160] = 16'hd0e5; data[161] = 16'h4efb; data[162] = 16'h4988; data[163] = 16'h0000;
	data[164] = 16'h0000; data[165] = 16'h0000; data[166] = 16'h0000; data[167] = 16'h0000;

	data[168] = 16'hd012; data[169] = 16'h5035; data[170] = 16'h4cad; data[171] = 16'h0000;
	data[172] = 16'h0000; data[173] = 16'h0000; data[174] = 16'h0000; data[175] = 16'h0000;
	data[176] = 16'hd05e; data[177] = 16'h4f76; data[178] = 16'h4bdc; data[179] = 16'h0000;
	data[180] = 16'h0000; data[181] = 16'h0000; data[182] = 16'h0000; data[183] = 16'h0000;
	data[184] = 16'hcfee; data[185] = 16'h4ffd; data[186] = 16'h4b86; data[187] = 16'h0000;
	data[188] = 16'h0000; data[189] = 16'h0000; data[190] = 16'h0000; data[191] = 16'h0000;

	data[192] = 16'hd041; data[193] = 16'h4ff3; data[194] = 16'h4c36; data[195] = 16'h0000;
	data[196] = 16'h0000; data[197] = 16'h0000; data[198] = 16'h0000; data[199] = 16'h0000;
	data[200] = 16'hd11b; data[201] = 16'h4de2; data[202] = 16'h48c0; data[203] = 16'h0000;
	data[204] = 16'h0000; data[205] = 16'h0000; data[206] = 16'h0000; data[207] = 16'h0000;
	data[208] = 16'hd1a2; data[209] = 16'h4c5c; data[210] = 16'h4237; data[211] = 16'h0000;
	data[212] = 16'h0000; data[213] = 16'h0000; data[214] = 16'h0000; data[215] = 16'h0000;

	weight[0] = 16'h341E; weight[1] = 16'h3867; weight[2] = 16'h3509; weight[3] = 16'h0000;
	weight[4] = 16'h0000; weight[5] = 16'h0000; weight[6] = 16'h0000; weight[7] = 16'h0000;
	weight[8] = 16'hAE6E; weight[9] = 16'hB0BF;	weight[10] = 16'hB0F7; weight[11] = 16'h0000;
	weight[12] = 16'h0000; weight[13] = 16'h0000; weight[14] = 16'h0000; weight[15] = 16'h0000;
	weight[16] = 16'hAC84; weight[17] = 16'hB2B4; weight[18] = 16'hAF54; weight[19] = 16'h0000;
	weight[20] = 16'h0000; weight[21] = 16'h0000; weight[22] = 16'h0000; weight[23] = 16'h0000;

	weight[24] = 16'h35C0; weight[25] = 16'h396D; weight[26] = 16'h36E1; weight[27] = 16'h0000;
	weight[28] = 16'h0000; weight[29] = 16'h0000; weight[30] = 16'h0000; weight[31] = 16'h0000;
	weight[32] = 16'hB10F; weight[33] = 16'hB456; weight[34] = 16'hB2C4; weight[35] = 16'h0000;
	weight[36] = 16'h0000; weight[37] = 16'h0000; weight[38] = 16'h0000; weight[39] = 16'h0000;
	weight[40] = 16'hB209; weight[41] = 16'hB76D; weight[42] = 16'hB3F0; weight[43] = 16'h0000;
	weight[44] = 16'h0000; weight[45] = 16'h0000; weight[46] = 16'h0000; weight[47] = 16'h0000;

	weight[48] = 16'h3282; weight[49] = 16'h376F; weight[50] = 16'h3504; weight[51] = 16'h0000;
	weight[52] = 16'h0000; weight[53] = 16'h0000; weight[54] = 16'h0000; weight[55] = 16'h0000;
	weight[56] = 16'hAE46; weight[57] = 16'hB1E7; weight[58] = 16'hACF0; weight[59] = 16'h0000;
	weight[60] = 16'h0000; weight[61] = 16'h0000; weight[62] = 16'h0000; weight[63] = 16'h0000;
	weight[64] = 16'hB249; weight[65] = 16'hB72B; weight[66] = 16'hB338; weight[67] = 16'h0000;
	weight[68] = 16'h0000; weight[69] = 16'h0000; weight[70] = 16'h0000; weight[71] = 16'h0000;*/
	data[0] = 16'h0000; data[1] = 16'h0000; data[2] = 16'h0000; data[3] = 16'h0000; data[4] = 16'h0000; data[5] = 16'h0000; data[6] = 16'h0000; data[7] = 16'h0000; data[8] = 16'h0000; data[9] = 16'h0000; data[10] = 16'h0000; data[11] = 16'h0000; data[12] = 16'h0000; data[13] = 16'h0000; data[14] = 16'h0000; data[15] = 16'h0000; data[16] = 16'h0000; data[17] = 16'h0000; data[18] = 16'h0000; data[19] = 16'h0000; data[20] = 16'h0000; data[21] = 16'h0000; data[22] = 16'h0000; data[23] = 16'h0000; data[24] = 16'h0000; data[25] = 16'h0000; data[26] = 16'h0000; data[27] = 16'h0000; data[28] = 16'h0000; data[29] = 16'h0000; data[30] = 16'h0000; data[31] = 16'h0000; data[32] = 16'h4dd3; data[33] = 16'h0000; data[34] = 16'h0000; data[35] = 16'h50b8; data[36] = 16'h55c6; data[37] = 16'h4c84; data[38] = 16'h5dee; data[39] = 16'h5593; data[40] = 16'h4e5b; data[41] = 16'h4c1f; data[42] = 16'h0000; data[43] = 16'h3c74; data[44] = 16'h566c; data[45] = 16'h4c65; data[46] = 16'h5e07; data[47] = 16'h50c1; data[48] = 16'h0000; data[49] = 16'h0000; data[50] = 16'h0000; data[51] = 16'h0000; data[52] = 16'h0000; data[53] = 16'h0000; data[54] = 16'h0000; data[55] = 16'h0000; data[56] = 16'h0000; data[57] = 16'h0000; data[58] = 16'h0000; data[59] = 16'h5238; data[60] = 16'h59fe; data[61] = 16'h4a36; data[62] = 16'h5d9c; data[63] = 16'h5acf; data[64] = 16'h0000; data[65] = 16'h0000; data[66] = 16'h0000; data[67] = 16'h0000; data[68] = 16'h5a43; data[69] = 16'h0000; data[70] = 16'h5db7; data[71] = 16'h5b44; data[72] = 16'h0000; data[73] = 16'h0000; data[74] = 16'h0000; data[75] = 16'h0000; data[76] = 16'h0000; data[77] = 16'h0000; data[78] = 16'h0000; data[79] = 16'h0000; data[80] = 16'h54ed; data[81] = 16'h0000; data[82] = 16'h0000; data[83] = 16'h5418; data[84] = 16'h5a51; data[85] = 16'h4cc1; data[86] = 16'h5da0; data[87] = 16'h5868; data[88] = 16'h54b9; data[89] = 16'h0000; data[90] = 16'h0000; data[91] = 16'h0000; data[92] = 16'h5a8e; data[93] = 16'h4a6e; data[94] = 16'h5d6f; data[95] = 16'h5a11; data[96] = 16'h0000; data[97] = 16'h0000; data[98] = 16'h0000; data[99] = 16'h0000; data[100] = 16'h0000; data[101] = 16'h0000; data[102] = 16'h0000; data[103] = 16'h0000; data[104] = 16'h5028; data[105] = 16'h0000; data[106]
= 16'h0000; data[107] = 16'h0000; data[108] = 16'h594c; data[109] = 16'h3bb8; data[110] = 16'h5da8; data[111] = 16'h5ade; data[112] = 16'h51d2;
data[113] = 16'h5001; data[114] = 16'h0000; data[115] = 16'h0000; data[116] = 16'h582c; data[117] = 16'h0000; data[118] = 16'h5d4d; data[119] =
16'h58b0; data[120] = 16'h0000; data[121] = 16'h0000; data[122] = 16'h0000; data[123] = 16'h0000; data[124] = 16'h0000; data[125] = 16'h0000; data[126] = 16'h0000; data[127] = 16'h0000; data[128] = 16'h0000; data[129] = 16'h48a3; data[130] = 16'h0000; data[131] = 16'h0000; data[132] = 16'h590c; data[133] = 16'h4c37; data[134] = 16'h5d01; data[135] = 16'h58cc; data[136] = 16'h5470; data[137] = 16'h5508; data[138] = 16'h0000; data[139] = 16'h0000; data[140] = 16'h5888; data[141] = 16'h4d39; data[142]
= 16'h5d48; data[143] = 16'h55d7; data[144] = 16'h0000; data[145] = 16'h0000; data[146] = 16'h0000; data[147] = 16'h0000; data[148] = 16'h0000;
data[149] = 16'h0000; data[150] = 16'h0000; data[151] = 16'h0000; data[152] = 16'h458c; data[153] = 16'h0000; data[154] = 16'h0000; data[155] =
16'h0000; data[156] = 16'h587a; data[157] = 16'h46fa; data[158] = 16'h5d2b; data[159] = 16'h5825; data[160] = 16'h5457; data[161] = 16'h55cc; data[162] = 16'h0000; data[163] = 16'h0000; data[164] = 16'h58d7; data[165] = 16'h5040; data[166] = 16'h5e1d; data[167] = 16'h552a; data[168] = 16'h0000; data[169] = 16'h0000; data[170] = 16'h0000; data[171] = 16'h0000; data[172] = 16'h0000; data[173] = 16'h0000; data[174] = 16'h0000; data[175] = 16'h0000; data[176] = 16'h5190; data[177] = 16'h0000; data[178]
= 16'h0000; data[179] = 16'h4c91; data[180] = 16'h56b9; data[181] = 16'h4e94; data[182] = 16'h5c27; data[183] = 16'h548a; data[184] = 16'h4ea3;
data[185] = 16'h53fb; data[186] = 16'h0000; data[187] = 16'h0000; data[188] = 16'h550d; data[189] = 16'h4f8e; data[190] = 16'h5d06; data[191] =
16'h542f; data[192] = 16'h0000; data[193] = 16'h0000; data[194] = 16'h0000; data[195] = 16'h0000; data[196] = 16'h0000; data[197] = 16'h0000; data[198] = 16'h0000; data[199] = 16'h0000; data[200] = 16'h56cb; data[201] = 16'h0000; data[202] = 16'h0000; data[203] = 16'h5093; data[204] = 16'h583f; data[205] = 16'h520b; data[206] = 16'h5c87; data[207] = 16'h5246; data[208] = 16'h5538; data[209] = 16'h0000; data[210] = 16'h0000; data[211] = 16'h0000; data[212] = 16'h575b; data[213] = 16'h5089; data[214]
= 16'h5cf5; data[215] = 16'h5374; data[216] = 16'h0000; data[217] = 16'h0000; data[218] = 16'h0000; data[219] = 16'h0000; data[220] = 16'h0000;
data[221] = 16'h0000; data[222] = 16'h0000; data[223] = 16'h0000; data[224] = 16'h53b0; data[225] = 16'h0000; data[226] = 16'h0000; data[227] =
16'h0000; data[228] = 16'h5431; data[229] = 16'h5110; data[230] = 16'h5e20; data[231] = 16'h533c; data[232] = 16'h537a; data[233] = 16'h0000; data[234] = 16'h0000; data[235] = 16'h0000; data[236] = 16'h580c; data[237] = 16'h0000; data[238] = 16'h5d27; data[239] = 16'h552c; data[240] = 16'h0000; data[241] = 16'h0000; data[242] = 16'h0000; data[243] = 16'h0000; data[244] = 16'h0000; data[245] = 16'h0000; data[246] = 16'h0000; data[247] = 16'h0000; data[248] = 16'h59b8; data[249] = 16'h0000; data[250]
= 16'h0000; data[251] = 16'h0000; data[252] = 16'h5914; data[253] = 16'h0000; data[254] = 16'h5ea3; data[255] = 16'h46bc; data[256] = 16'h580f;
data[257] = 16'h0000; data[258] = 16'h0000; data[259] = 16'h0000; data[260] = 16'h564c; data[261] = 16'h0000; data[262] = 16'h5d4e; data[263] =
16'h4c00; data[264] = 16'h0000; data[265] = 16'h0000; data[266] = 16'h0000; data[267] = 16'h0000; data[268] = 16'h0000; data[269] = 16'h0000; data[270] = 16'h0000; data[271] = 16'h0000; data[272] = 16'h5b79; data[273] = 16'h0000; data[274] = 16'h0000; data[275] = 16'h0000; data[276] = 16'h596d; data[277] = 16'h4aa2; data[278] = 16'h5c94; data[279] = 16'h0000; data[280] = 16'h5827; data[281] = 16'h0000; data[282] = 16'h0000; data[283] = 16'h0000; data[284] = 16'h566d; data[285] = 16'h492b; data[286]
= 16'h5d45; data[287] = 16'h4fd2; data[288] = 16'h0000; data[289] = 16'h0000; data[290] = 16'h0000; data[291] = 16'h0000; data[292] = 16'h0000;
data[293] = 16'h0000; data[294] = 16'h0000; data[295] = 16'h0000; data[296] = 16'h5713; data[297] = 16'h0000; data[298] = 16'h0000; data[299] =
16'h579f; data[300] = 16'h55ac; data[301] = 16'h5164; data[302] = 16'h5cf8; data[303] = 16'h512a; data[304] = 16'h5763; data[305] = 16'h0000; data[306] = 16'h0000; data[307] = 16'h0000; data[308] = 16'h562b; data[309] = 16'h500a; data[310] = 16'h5c71; data[311] = 16'h51dd; data[312] = 16'h0000; data[313] = 16'h0000; data[314] = 16'h0000; data[315] = 16'h0000; data[316] = 16'h0000; data[317] = 16'h0000; data[318] = 16'h0000; data[319] = 16'h0000; data[320] = 16'h5147; data[321] = 16'h0000; data[322]
= 16'h49db; data[323] = 16'h5613; data[324] = 16'h5545; data[325] = 16'h5145; data[326] = 16'h5ce2; data[327] = 16'h564b; data[328] = 16'h4f72;
data[329] = 16'h0000; data[330] = 16'h0000; data[331] = 16'h4df8; data[332] = 16'h54ee; data[333] = 16'h52c6; data[334] = 16'h5cba; data[335] =
16'h5504; data[336] = 16'h0000; data[337] = 16'h0000; data[338] = 16'h0000; data[339] = 16'h0000; data[340] = 16'h0000; data[341] = 16'h0000; data[342] = 16'h0000; data[343] = 16'h0000; data[344] = 16'h45c8; data[345] = 16'h0000; data[346] = 16'h47d7; data[347] = 16'h4cd3; data[348] = 16'h5415; data[349] = 16'h50d4; data[350] = 16'h5cd8; data[351] = 16'h57e3; data[352] = 16'h5348; data[353] = 16'h0000; data[354] = 16'h0000; data[355] = 16'h0000; data[356] = 16'h5621; data[357] = 16'h4baf; data[358]
= 16'h5d0b; data[359] = 16'h5390; data[360] = 16'h0000; data[361] = 16'h0000; data[362] = 16'h0000; data[363] = 16'h0000; data[364] = 16'h0000;
data[365] = 16'h0000; data[366] = 16'h0000; data[367] = 16'h0000; data[368] = 16'h4f8e; data[369] = 16'h0000; data[370] = 16'h0000; data[371] =
16'h482e; data[372] = 16'h54b8; data[373] = 16'h499b; data[374] = 16'h5cb8; data[375] = 16'h54b2; data[376] = 16'h5460; data[377] = 16'h0000; data[378] = 16'h0000; data[379] = 16'h0000; data[380] = 16'h55e5; data[381] = 16'h470f; data[382] = 16'h5cb6; data[383] = 16'h5498; data[384] = 16'h0000; data[385] = 16'h0000; data[386] = 16'h0000; data[387] = 16'h0000; data[388] = 16'h0000; data[389] = 16'h0000; data[390] = 16'h0000; data[391] = 16'h0000; data[392] = 16'h50e7; data[393] = 16'h40c4; data[394]
= 16'h0000; data[395] = 16'h0000; data[396] = 16'h5539; data[397] = 16'h507a; data[398] = 16'h5d37; data[399] = 16'h512b; data[400] = 16'h5347;
data[401] = 16'h5012; data[402] = 16'h0000; data[403] = 16'h0000; data[404] = 16'h55f4; data[405] = 16'h4c0f; data[406] = 16'h5d6f; data[407] =
16'h5397; data[408] = 16'h0000; data[409] = 16'h0000; data[410] = 16'h0000; data[411] = 16'h0000; data[412] = 16'h0000; data[413] = 16'h0000; data[414] = 16'h0000; data[415] = 16'h0000; data[416] = 16'h4f41; data[417] = 16'h4bea; data[418] = 16'h4d21; data[419] = 16'h0000; data[420] = 16'h529d; data[421] = 16'h50b2; data[422] = 16'h5d58; data[423] = 16'h54f0; data[424] = 16'h54ac; data[425] = 16'h5699; data[426] = 16'h0000; data[427] = 16'h0000; data[428] = 16'h584e; data[429] = 16'h0000; data[430]
= 16'h5db7; data[431] = 16'h534a; data[432] = 16'h0000; data[433] = 16'h0000; data[434] = 16'h0000; data[435] = 16'h0000; data[436] = 16'h0000;
data[437] = 16'h0000; data[438] = 16'h0000; data[439] = 16'h0000; data[440] = 16'h4f86; data[441] = 16'h0000; data[442] = 16'h49b9; data[443] =
16'h0000; data[444] = 16'h54f2; data[445] = 16'h4bd8; data[446] = 16'h5d21; data[447] = 16'h56ec; data[448] = 16'h57fc; data[449] = 16'h5605; data[450] = 16'h0000; data[451] = 16'h0000; data[452] = 16'h5c8a; data[453] = 16'h4b94; data[454] = 16'h5d27; data[455] = 16'h5510; data[456] = 16'h0000; data[457] = 16'h0000; data[458] = 16'h0000; data[459] = 16'h0000; data[460] = 16'h0000; data[461] = 16'h0000; data[462] = 16'h0000; data[463] = 16'h0000; data[464] = 16'h5634; data[465] = 16'h0000; data[466]
= 16'h0000; data[467] = 16'h0000; data[468] = 16'h5807; data[469] = 16'h50e3; data[470] = 16'h5cf6; data[471] = 16'h5598; data[472] = 16'h5664;
data[473] = 16'h48d0; data[474] = 16'h0000; data[475] = 16'h0000; data[476] = 16'h5cba; data[477] = 16'h4c28; data[478] = 16'h5cf3; data[479] =
16'h58a9; data[480] = 16'h0000; data[481] = 16'h0000; data[482] = 16'h0000; data[483] = 16'h0000; data[484] = 16'h0000; data[485] = 16'h0000; data[486] = 16'h0000; data[487] = 16'h0000; data[488] = 16'h55a0; data[489] = 16'h0000; data[490] = 16'h0000; data[491] = 16'h0000; data[492] = 16'h5807; data[493] = 16'h4fbc; data[494] = 16'h5dad; data[495] = 16'h55db; data[496] = 16'h5686; data[497] = 16'h0000; data[498] = 16'h0000; data[499] = 16'h0000; data[500] = 16'h58cc; data[501] = 16'h5057; data[502]
= 16'h5dbc; data[503] = 16'h557f; data[504] = 16'h0000; data[505] = 16'h0000; data[506] = 16'h0000; data[507] = 16'h0000; data[508] = 16'h0000;
data[509] = 16'h0000; data[510] = 16'h0000; data[511] = 16'h0000; data[512] = 16'h4f16; data[513] = 16'h0000; data[514] = 16'h0000; data[515] =
16'h0000; data[516] = 16'h5615; data[517] = 16'h4b90; data[518] = 16'h5dbb; data[519] = 16'h55c7; data[520] = 16'h54a6; data[521] = 16'h0000; data[522] = 16'h0000; data[523] = 16'h4d49; data[524] = 16'h5622; data[525] = 16'h4d0e; data[526] = 16'h5d89; data[527] = 16'h53ac; data[528] = 16'h0000; data[529] = 16'h0000; data[530] = 16'h0000; data[531] = 16'h0000; data[532] = 16'h0000; data[533] = 16'h0000; data[534] = 16'h0000; data[535] = 16'h0000; data[536] = 16'h5064; data[537] = 16'h0000; data[538]
= 16'h0000; data[539] = 16'h0000; data[540] = 16'h5667; data[541] = 16'h4a17; data[542] = 16'h5ca1; data[543] = 16'h5531; data[544] = 16'h45ca;
data[545] = 16'h0000; data[546] = 16'h0000; data[547] = 16'h5012; data[548] = 16'h55bc; data[549] = 16'h4de2; data[550] = 16'h5d51; data[551] =
16'h5518; data[552] = 16'h0000; data[553] = 16'h0000; data[554] = 16'h0000; data[555] = 16'h0000; data[556] = 16'h0000; data[557] = 16'h0000; data[558] = 16'h0000; data[559] = 16'h0000; data[560] = 16'h572c; data[561] = 16'h0000; data[562] = 16'h0000; data[563] = 16'h0000; data[564] = 16'h5739; data[565] = 16'h4ad4; data[566] = 16'h5d75; data[567] = 16'h51bc; data[568] = 16'h53cd; data[569] = 16'h0000; data[570] = 16'h0000; data[571] = 16'h4d5a; data[572] = 16'h5665; data[573] = 16'h4c81; data[574]
= 16'h5de3; data[575] = 16'h5418; data[576] = 16'h0000; data[577] = 16'h0000; data[578] = 16'h0000; data[579] = 16'h0000; data[580] = 16'h0000;
data[581] = 16'h0000; data[582] = 16'h0000; data[583] = 16'h0000; data[584] = 16'h51e6; data[585] = 16'h0000; data[586] = 16'h0000; data[587] =
16'h0000; data[588] = 16'h57ad; data[589] = 16'h4d1e; data[590] = 16'h5d61; data[591] = 16'h55cf; data[592] = 16'h38c0; data[593] = 16'h0000; data[594] = 16'h0000; data[595] = 16'h0000; data[596] = 16'h5688; data[597] = 16'h49df; data[598] = 16'h5dd3; data[599] = 16'h579c; data[600] = 16'h0000; data[601] = 16'h0000; data[602] = 16'h0000; data[603] = 16'h0000; data[604] = 16'h0000; data[605] = 16'h0000; data[606] = 16'h0000; data[607] = 16'h0000; data[608] = 16'h4903; data[609] = 16'h4191; data[610]
= 16'h0000; data[611] = 16'h0000; data[612] = 16'h5487; data[613] = 16'h5019; data[614] = 16'h5d97; data[615] = 16'h5612; data[616] = 16'h0000;
data[617] = 16'h0000; data[618] = 16'h0000; data[619] = 16'h0000; data[620] = 16'h5512; data[621] = 16'h50bf; data[622] = 16'h5d3d; data[623] =
16'h5747; data[624] = 16'h0000; data[625] = 16'h0000; data[626] = 16'h0000; data[627] = 16'h0000; data[628] = 16'h0000; data[629] = 16'h0000; data[630] = 16'h0000; data[631] = 16'h0000; data[632] = 16'h54a4; data[633] = 16'h0000; data[634] = 16'h0000; data[635] = 16'h0000; data[636] = 16'h580d; data[637] = 16'h4bfe; data[638] = 16'h5d79; data[639] = 16'h5522; data[640] = 16'h5481; data[641] = 16'h0000; data[642] = 16'h0000; data[643] = 16'h0000; data[644] = 16'h5966; data[645] = 16'h4dac; data[646]
= 16'h5d30; data[647] = 16'h5546; data[648] = 16'h0000; data[649] = 16'h0000; data[650] = 16'h0000; data[651] = 16'h0000; data[652] = 16'h0000;
data[653] = 16'h0000; data[654] = 16'h0000; data[655] = 16'h0000; data[656] = 16'h52d7; data[657] = 16'h0000; data[658] = 16'h0000; data[659] =
16'h0000; data[660] = 16'h5652; data[661] = 16'h50d9; data[662] = 16'h5cac; data[663] = 16'h54e8; data[664] = 16'h5565; data[665] = 16'h0000; data[666] = 16'h0000; data[667] = 16'h0000; data[668] = 16'h58cf; data[669] = 16'h4cf5; data[670] = 16'h5d37; data[671] = 16'h5384; data[672] = 16'h0000; data[673] = 16'h0000; data[674] = 16'h0000; data[675] = 16'h0000; data[676] = 16'h0000; data[677] = 16'h0000; data[678] = 16'h0000; data[679] = 16'h0000; data[680] = 16'h5307; data[681] = 16'h0000; data[682]
= 16'h48de; data[683] = 16'h4d00; data[684] = 16'h51d0; data[685] = 16'h5044; data[686] = 16'h5d6f; data[687] = 16'h5253; data[688] = 16'h5128;
data[689] = 16'h0000; data[690] = 16'h0000; data[691] = 16'h55d4; data[692] = 16'h561e; data[693] = 16'h46a0; data[694] = 16'h5e30; data[695] =
16'h5a31; data[696] = 16'h0000; data[697] = 16'h0000; data[698] = 16'h0000; data[699] = 16'h0000; data[700] = 16'h0000; data[701] = 16'h0000; data[702] = 16'h0000; data[703] = 16'h0000; data[704] = 16'h4e3f; data[705] = 16'h0000; data[706] = 16'h4f53; data[707] = 16'h52d0; data[708] = 16'h51b7; data[709] = 16'h4d7e; data[710] = 16'h5dcf; data[711] = 16'h5610; data[712] = 16'h0000; data[713] = 16'h0000; data[714] = 16'h55d3; data[715] = 16'h5a84; data[716] = 16'h5530; data[717] = 16'h5422; data[718]
= 16'h5e1c; data[719] = 16'h5c53; data[720] = 16'h0000; data[721] = 16'h0000; data[722] = 16'h0000; data[723] = 16'h0000; data[724] = 16'h0000;
data[725] = 16'h0000; data[726] = 16'h0000; data[727] = 16'h0000; data[728] = 16'h0000; data[729] = 16'h0000; data[730] = 16'h5293; data[731] =
16'h58f7; data[732] = 16'h562f; data[733] = 16'h4f5a; data[734] = 16'h5ddb; data[735] = 16'h5bb9; data[736] = 16'h0000; data[737] = 16'h0000; data[738] = 16'h55a9; data[739] = 16'h5ad0; data[740] = 16'h55f4; data[741] = 16'h554c; data[742] = 16'h5c1f; data[743] = 16'h5c42; data[744] = 16'h0000; data[745] = 16'h0000; data[746] = 16'h0000; data[747] = 16'h0000; data[748] = 16'h0000; data[749] = 16'h0000; data[750] = 16'h0000; data[751] = 16'h0000; data[752] = 16'h50dc; data[753] = 16'h0000; data[754]
= 16'h54f3; data[755] = 16'h59de; data[756] = 16'h5608; data[757] = 16'h54ea; data[758] = 16'h5c9e; data[759] = 16'h59a1; data[760] = 16'h0000;
data[761] = 16'h0000; data[762] = 16'h5419; data[763] = 16'h5935; data[764] = 16'h5597; data[765] = 16'h5404; data[766] = 16'h550a; data[767] =
16'h5b59; data[768] = 16'h0000; data[769] = 16'h0000; data[770] = 16'h0000; data[771] = 16'h0000; data[772] = 16'h0000; data[773] = 16'h0000; data[774] = 16'h0000; data[775] = 16'h0000; data[776] = 16'h5a8b; data[777] = 16'h0000; data[778] = 16'h58e9; data[779] = 16'h5a02; data[780] = 16'h5464; data[781] = 16'h586d; data[782] = 16'h5bb5; data[783] = 16'h4e8b; data[784] = 16'h5863; data[785] = 16'h0000; data[786] = 16'h582a; data[787] = 16'h560f; data[788] = 16'h50a4; data[789] = 16'h5810; data[790]
= 16'h52b2; data[791] = 16'h4cd7; data[792] = 16'h0000; data[793] = 16'h0000; data[794] = 16'h0000; data[795] = 16'h0000; data[796] = 16'h0000;
data[797] = 16'h0000; data[798] = 16'h0000; data[799] = 16'h0000; data[800] = 16'h5c99; data[801] = 16'h0000; data[802] = 16'h5431; data[803] =
16'h5aa7; data[804] = 16'h55c0; data[805] = 16'h56b3; data[806] = 16'h5ced; data[807] = 16'h0000; data[808] = 16'h5bc7; data[809] = 16'h0000; data[810] = 16'h566d; data[811] = 16'h5a81; data[812] = 16'h56f6; data[813] = 16'h5844; data[814] = 16'h5703; data[815] = 16'h0000; data[816] = 16'h0000; data[817] = 16'h0000; data[818] = 16'h0000; data[819] = 16'h0000; data[820] = 16'h0000; data[821] = 16'h0000; data[822] = 16'h0000; data[823] = 16'h0000; data[824] = 16'h5795; data[825] = 16'h0000; data[826]
= 16'h5126; data[827] = 16'h5565; data[828] = 16'h5564; data[829] = 16'h53e0; data[830] = 16'h5cd4; data[831] = 16'h50fc; data[832] = 16'h5c85;
data[833] = 16'h0000; data[834] = 16'h4f55; data[835] = 16'h5bb9; data[836] = 16'h5875; data[837] = 16'h58b8; data[838] = 16'h59c4; data[839] =
16'h0000; data[840] = 16'h0000; data[841] = 16'h0000; data[842] = 16'h0000; data[843] = 16'h0000; data[844] = 16'h0000; data[845] = 16'h0000; data[846] = 16'h0000; data[847] = 16'h0000; data[848] = 16'h5796; data[849] = 16'h0000; data[850] = 16'h0000; data[851] = 16'h5047; data[852] = 16'h5547; data[853] = 16'h537d; data[854] = 16'h5cdd; data[855] = 16'h3f5c; data[856] = 16'h5daf; data[857] = 16'h0000; data[858] = 16'h0000; data[859] = 16'h5b8f; data[860] = 16'h590c; data[861] = 16'h580c; data[862]
= 16'h5c21; data[863] = 16'h0000; data[864] = 16'h0000; data[865] = 16'h0000; data[866] = 16'h0000; data[867] = 16'h0000; data[868] = 16'h0000;
data[869] = 16'h0000; data[870] = 16'h0000; data[871] = 16'h0000; data[872] = 16'h5426; data[873] = 16'h0000; data[874] = 16'h0000; data[875] =
16'h4ef4; data[876] = 16'h56d5; data[877] = 16'h5076; data[878] = 16'h5c46; data[879] = 16'h50c2; data[880] = 16'h5715; data[881] = 16'h0000; data[882] = 16'h0000; data[883] = 16'h5394; data[884] = 16'h56c3; data[885] = 16'h53b1; data[886] = 16'h5bad; data[887] = 16'h4e12; data[888] = 16'h0000; data[889] = 16'h0000; data[890] = 16'h0000; data[891] = 16'h0000; data[892] = 16'h0000; data[893] = 16'h0000; data[894] = 16'h0000; data[895] = 16'h0000; data[896] = 16'h5540; data[897] = 16'h0000; data[898]
= 16'h0000; data[899] = 16'h4fac; data[900] = 16'h55b0; data[901] = 16'h5056; data[902] = 16'h5c0f; data[903] = 16'h4fc3; data[904] = 16'h5204;
data[905] = 16'h0000; data[906] = 16'h0000; data[907] = 16'h4b3c; data[908] = 16'h5800; data[909] = 16'h4f63; data[910] = 16'h5a92; data[911] =
16'h5378; data[912] = 16'h0000; data[913] = 16'h0000; data[914] = 16'h0000; data[915] = 16'h0000; data[916] = 16'h0000; data[917] = 16'h0000; data[918] = 16'h0000; data[919] = 16'h0000; data[920] = 16'h5155; data[921] = 16'h0000; data[922] = 16'h0000; data[923] = 16'h4d33; data[924] = 16'h5525; data[925] = 16'h4e59; data[926] = 16'h5b0a; data[927] = 16'h5497; data[928] = 16'h52b8; data[929] = 16'h0000; data[930] = 16'h0000; data[931] = 16'h4d56; data[932] = 16'h5504; data[933] = 16'h4cc2; data[934]
= 16'h5ae1; data[935] = 16'h52dc; data[936] = 16'h0000; data[937] = 16'h0000; data[938] = 16'h0000; data[939] = 16'h0000; data[940] = 16'h0000;
data[941] = 16'h0000; data[942] = 16'h0000; data[943] = 16'h0000; data[944] = 16'h5291; data[945] = 16'h0000; data[946] = 16'h4b64; data[947] =
16'h4d42; data[948] = 16'h530e; data[949] = 16'h5085; data[950] = 16'h5ba6; data[951] = 16'h5390; data[952] = 16'h5210; data[953] = 16'h3960; data[954] = 16'h0000; data[955] = 16'h4734; data[956] = 16'h55b7; data[957] = 16'h4e93; data[958] = 16'h5a93; data[959] = 16'h5507; data[960] = 16'h0000; data[961] = 16'h0000; data[962] = 16'h0000; data[963] = 16'h0000; data[964] = 16'h0000; data[965] = 16'h0000; data[966] = 16'h0000; data[967] = 16'h0000; data[968] = 16'h526e; data[969] = 16'h4cf0; data[970]
= 16'h0000; data[971] = 16'h0000; data[972] = 16'h52fe; data[973] = 16'h4e4d; data[974] = 16'h5bbc; data[975] = 16'h5068; data[976] = 16'h5093;
data[977] = 16'h0000; data[978] = 16'h0000; data[979] = 16'h5198; data[980] = 16'h55dc; data[981] = 16'h4fc0; data[982] = 16'h5bab; data[983] =
16'h5542; data[984] = 16'h0000; data[985] = 16'h0000; data[986] = 16'h0000; data[987] = 16'h0000; data[988] = 16'h0000; data[989] = 16'h0000; data[990] = 16'h0000; data[991] = 16'h0000; data[992] = 16'h5334; data[993] = 16'h0000; data[994] = 16'h4069; data[995] = 16'h31b0; data[996] = 16'h5072; data[997] = 16'h4c8a; data[998] = 16'h5bee; data[999] = 16'h4c3f; data[1000] = 16'h51fb; data[1001] = 16'h0000; data[1002] = 16'h0000; data[1003] = 16'h504b; data[1004] = 16'h51df; data[1005] = 16'h4d25; data[1006] = 16'h5be2; data[1007] = 16'h4dbe; data[1008] = 16'h0000; data[1009] = 16'h0000; data[1010] = 16'h0000; data[1011] = 16'h0000; data[1012] = 16'h0000; data[1013] = 16'h0000; data[1014] = 16'h0000; data[1015] =
16'h0000; data[1016] = 16'h5505; data[1017] = 16'h0000; data[1018] = 16'h405b; data[1019] = 16'h4ca2; data[1020] = 16'h5339; data[1021] = 16'h4cca; data[1022] = 16'h5b80; data[1023] = 16'h4d71; data[1024] = 16'h4f0b; data[1025] = 16'h5141; data[1026] = 16'h0000; data[1027] = 16'h0000; data[1028] = 16'h530d; data[1029] = 16'h4fc3; data[1030] = 16'h5b5b; data[1031] = 16'h51c2; data[1032] = 16'h0000; data[1033] = 16'h0000; data[1034] = 16'h0000; data[1035] = 16'h0000; data[1036] = 16'h0000; data[1037]
= 16'h0000; data[1038] = 16'h0000; data[1039] = 16'h0000; data[1040] = 16'h51a4; data[1041] = 16'h0000; data[1042] = 16'h0000; data[1043] = 16'h0000; data[1044] = 16'h54fa; data[1045] = 16'h4e25; data[1046] = 16'h5b32; data[1047] = 16'h5558; data[1048] = 16'h50dc; data[1049] = 16'h5287;
data[1050] = 16'h4bc0; data[1051] = 16'h0000; data[1052] = 16'h51c6; data[1053] = 16'h5041; data[1054] = 16'h5bef; data[1055] = 16'h53c9; data[1056] = 16'h0000; data[1057] = 16'h0000; data[1058] = 16'h0000; data[1059] = 16'h0000; data[1060] = 16'h0000; data[1061] = 16'h0000; data[1062] = 16'h0000; data[1063] = 16'h0000; data[1064] = 16'h5450; data[1065] = 16'h0000; data[1066] = 16'h0000; data[1067] = 16'h4f04; data[1068] = 16'h5418; data[1069] = 16'h4e7a; data[1070] = 16'h5c1f; data[1071] = 16'h5120; data[1072] = 16'h5418; data[1073] = 16'h0000; data[1074] = 16'h0000; data[1075] = 16'h4718; data[1076] = 16'h5354; data[1077] = 16'h4c9e; data[1078] = 16'h5c02; data[1079] = 16'h4f22; data[1080] = 16'h0000; data[1081] = 16'h0000; data[1082] = 16'h0000; data[1083] = 16'h0000; data[1084] = 16'h0000; data[1085] = 16'h0000; data[1086] = 16'h0000; data[1087] =
16'h0000; data[1088] = 16'h50f2; data[1089] = 16'h0000; data[1090] = 16'h49a0; data[1091] = 16'h4d6c; data[1092] = 16'h521f; data[1093] = 16'h4cee; data[1094] = 16'h5c3b; data[1095] = 16'h5461; data[1096] = 16'h5392; data[1097] = 16'h0000; data[1098] = 16'h0000; data[1099] = 16'h0000; data[1100] = 16'h5328; data[1101] = 16'h4cf8; data[1102] = 16'h5a9a; data[1103] = 16'h5097; data[1104] = 16'h0000; data[1105] = 16'h0000; data[1106] = 16'h0000; data[1107] = 16'h0000; data[1108] = 16'h0000; data[1109]
= 16'h0000; data[1110] = 16'h0000; data[1111] = 16'h0000; data[1112] = 16'h4f34; data[1113] = 16'h0000; data[1114] = 16'h0000; data[1115] = 16'h4af4; data[1116] = 16'h55c2; data[1117] = 16'h4f83; data[1118] = 16'h5b65; data[1119] = 16'h56ac; data[1120] = 16'h5218; data[1121] = 16'h5046;
data[1122] = 16'h0000; data[1123] = 16'h0000; data[1124] = 16'h5584; data[1125] = 16'h4de7; data[1126] = 16'h5a07; data[1127] = 16'h5290; data[1128] = 16'h0000; data[1129] = 16'h0000; data[1130] = 16'h0000; data[1131] = 16'h0000; data[1132] = 16'h0000; data[1133] = 16'h0000; data[1134] = 16'h0000; data[1135] = 16'h0000; data[1136] = 16'h5314; data[1137] = 16'h521d; data[1138] = 16'h4c6f; data[1139] = 16'h0000; data[1140] = 16'h5290; data[1141] = 16'h505e; data[1142] = 16'h5c42; data[1143] = 16'h518a; data[1144] = 16'h517e; data[1145] = 16'h0000; data[1146] = 16'h0000; data[1147] = 16'h4f98; data[1148] = 16'h55d4; data[1149] = 16'h50d9; data[1150] = 16'h5c17; data[1151] = 16'h5612; data[1152] = 16'h0000; data[1153] = 16'h0000; data[1154] = 16'h0000; data[1155] = 16'h0000; data[1156] = 16'h0000; data[1157] = 16'h0000; data[1158] = 16'h0000; data[1159] =
16'h0000; data[1160] = 16'h5209; data[1161] = 16'h52e5; data[1162] = 16'h498e; data[1163] = 16'h0000; data[1164] = 16'h5268; data[1165] = 16'h4d20; data[1166] = 16'h5c84; data[1167] = 16'h50af; data[1168] = 16'h52a4; data[1169] = 16'h0000; data[1170] = 16'h0000; data[1171] = 16'h4e78; data[1172] = 16'h549c; data[1173] = 16'h4c02; data[1174] = 16'h5c93; data[1175] = 16'h54e8; data[1176] = 16'h0000; data[1177] = 16'h0000; data[1178] = 16'h0000; data[1179] = 16'h0000; data[1180] = 16'h0000; data[1181]
= 16'h0000; data[1182] = 16'h0000; data[1183] = 16'h0000; data[1184] = 16'h525c; data[1185] = 16'h5461; data[1186] = 16'h4096; data[1187] = 16'h0000; data[1188] = 16'h5377; data[1189] = 16'h4f89; data[1190] = 16'h5c6f; data[1191] = 16'h52c9; data[1192] = 16'h5072; data[1193] = 16'h4917;
data[1194] = 16'h0000; data[1195] = 16'h0000; data[1196] = 16'h53ca; data[1197] = 16'h4c29; data[1198] = 16'h5c6c; data[1199] = 16'h52ff; data[1200] = 16'h0000; data[1201] = 16'h0000; data[1202] = 16'h0000; data[1203] = 16'h0000; data[1204] = 16'h0000; data[1205] = 16'h0000; data[1206] = 16'h0000; data[1207] = 16'h0000; data[1208] = 16'h4e4c; data[1209] = 16'h4a90; data[1210] = 16'h4d6e; data[1211] = 16'h0000; data[1212] = 16'h53d4; data[1213] = 16'h532a; data[1214] = 16'h5d13; data[1215] = 16'h54f6; data[1216] = 16'h50f4; data[1217] = 16'h0000; data[1218] = 16'h476d; data[1219] = 16'h49eb; data[1220] = 16'h5193; data[1221] = 16'h50ba; data[1222] = 16'h5c7c; data[1223] = 16'h50eb; data[1224] = 16'h0000; data[1225] = 16'h0000; data[1226] = 16'h0000; data[1227] = 16'h0000; data[1228] = 16'h0000; data[1229] = 16'h0000; data[1230] = 16'h0000; data[1231] =
16'h0000; data[1232] = 16'h5280; data[1233] = 16'h5029; data[1234] = 16'h4880; data[1235] = 16'h0000; data[1236] = 16'h521d; data[1237] = 16'h4ff0; data[1238] = 16'h5d2f; data[1239] = 16'h50a2; data[1240] = 16'h51ee; data[1241] = 16'h4e85; data[1242] = 16'h4224; data[1243] = 16'h4e2b; data[1244] = 16'h51b0; data[1245] = 16'h507a; data[1246] = 16'h5cbd; data[1247] = 16'h4fb5; data[1248] = 16'h0000; data[1249] = 16'h0000; data[1250] = 16'h0000; data[1251] = 16'h0000; data[1252] = 16'h0000; data[1253]
= 16'h0000; data[1254] = 16'h0000; data[1255] = 16'h0000; data[1256] = 16'h52d8; data[1257] = 16'h4a4b; data[1258] = 16'h50f3; data[1259] = 16'h448b; data[1260] = 16'h5023; data[1261] = 16'h4f18; data[1262] = 16'h5cb5; data[1263] = 16'h50c0; data[1264] = 16'h51b3; data[1265] = 16'h4b6d;
data[1266] = 16'h468a; data[1267] = 16'h4916; data[1268] = 16'h5248; data[1269] = 16'h4d62; data[1270] = 16'h5c86; data[1271] = 16'h51dc; data[1272] = 16'h0000; data[1273] = 16'h0000; data[1274] = 16'h0000; data[1275] = 16'h0000; data[1276] = 16'h0000; data[1277] = 16'h0000; data[1278] = 16'h0000; data[1279] = 16'h0000; data[1280] = 16'h545e; data[1281] = 16'h4d2a; data[1282] = 16'h4b6a; data[1283] = 16'h0000; data[1284] = 16'h52c2; data[1285] = 16'h4bda; data[1286] = 16'h5c6c; data[1287] = 16'h4fa4; data[1288] = 16'h522d; data[1289] = 16'h48f3; data[1290] = 16'h0000; data[1291] = 16'h435c; data[1292] = 16'h529b; data[1293] = 16'h4cda; data[1294] = 16'h5b62; data[1295] = 16'h5072; data[1296] = 16'h0000; data[1297] = 16'h0000; data[1298] = 16'h0000; data[1299] = 16'h0000; data[1300] = 16'h0000; data[1301] = 16'h0000; data[1302] = 16'h0000; data[1303] =
16'h0000; data[1304] = 16'h5534; data[1305] = 16'h50d6; data[1306] = 16'h0000; data[1307] = 16'h0000; data[1308] = 16'h5613; data[1309] = 16'h4e54; data[1310] = 16'h5b4d; data[1311] = 16'h520d; data[1312] = 16'h525f; data[1313] = 16'h55a7; data[1314] = 16'h0000; data[1315] = 16'h0000; data[1316] = 16'h5529; data[1317] = 16'h4f76; data[1318] = 16'h5bab; data[1319] = 16'h50e7; data[1320] = 16'h0000; data[1321] = 16'h0000; data[1322] = 16'h0000; data[1323] = 16'h0000; data[1324] = 16'h0000; data[1325]
= 16'h0000; data[1326] = 16'h0000; data[1327] = 16'h0000; data[1328] = 16'h5440; data[1329] = 16'h0000; data[1330] = 16'h0000; data[1331] = 16'h54b5; data[1332] = 16'h57b0; data[1333] = 16'h5430; data[1334] = 16'h5ca3; data[1335] = 16'h5529; data[1336] = 16'h4f1c; data[1337] = 16'h5388;
data[1338] = 16'h4d5c; data[1339] = 16'h49d9; data[1340] = 16'h5390; data[1341] = 16'h51ce; data[1342] = 16'h5b5e; data[1343] = 16'h525f; data[1344] = 16'h0000; data[1345] = 16'h0000; data[1346] = 16'h0000; data[1347] = 16'h0000; data[1348] = 16'h0000; data[1349] = 16'h0000; data[1350] = 16'h0000; data[1351] = 16'h0000; data[1352] = 16'h5076; data[1353] = 16'h0000; data[1354] = 16'h4c00; data[1355] = 16'h5555; data[1356] = 16'h539b; data[1357] = 16'h5160; data[1358] = 16'h5cd4; data[1359] = 16'h554e; data[1360] = 16'h5066; data[1361] = 16'h515c; data[1362] = 16'h5046; data[1363] = 16'h4e67; data[1364] = 16'h518d; data[1365] = 16'h518b; data[1366] = 16'h5a9c; data[1367] = 16'h519d; data[1368] = 16'h0000; data[1369] = 16'h0000; data[1370] = 16'h0000; data[1371] = 16'h0000; data[1372] = 16'h0000; data[1373] = 16'h0000; data[1374] = 16'h0000; data[1375] =
16'h0000; data[1376] = 16'h0000; data[1377] = 16'h0000; data[1378] = 16'h0000; data[1379] = 16'h0000; data[1380] = 16'h0000; data[1381] = 16'h0000; data[1382] = 16'h0000; data[1383] = 16'h0000; data[1384] = 16'h0000; data[1385] = 16'h0000; data[1386] = 16'h0000; data[1387] = 16'h0000; data[1388] = 16'h0000; data[1389] = 16'h0000; data[1390] = 16'h0000; data[1391] = 16'h0000; data[1392] = 16'h0000; data[1393] = 16'h0000; data[1394] = 16'h0000; data[1395] = 16'h0000; data[1396] = 16'h0000; data[1397]
= 16'h0000; data[1398] = 16'h0000; data[1399] = 16'h0000; data[1400] = 16'h0000; data[1401] = 16'h0000; data[1402] = 16'h0000; data[1403] = 16'h0000; data[1404] = 16'h0000; data[1405] = 16'h0000; data[1406] = 16'h0000; data[1407] = 16'h0000; data[1408] = 16'h0000; data[1409] = 16'h0000;
data[1410] = 16'h0000; data[1411] = 16'h0000; data[1412] = 16'h0000; data[1413] = 16'h0000; data[1414] = 16'h0000; data[1415] = 16'h0000; data[1416] = 16'h0000; data[1417] = 16'h0000; data[1418] = 16'h0000; data[1419] = 16'h0000; data[1420] = 16'h0000; data[1421] = 16'h0000; data[1422] = 16'h0000; data[1423] = 16'h0000; data[1424] = 16'h52ef; data[1425] = 16'h505a; data[1426] = 16'h5572; data[1427] = 16'h51a8; data[1428] = 16'h55f1; data[1429] = 16'h507f; data[1430] = 16'h0000; data[1431] = 16'h50d3; data[1432] = 16'h5111; data[1433] = 16'h4ccb; data[1434] = 16'h548d; data[1435] = 16'h5294; data[1436] = 16'h55cb; data[1437] = 16'h5058; data[1438] = 16'h4c46; data[1439] = 16'h4eea; data[1440] = 16'h0000; data[1441] = 16'h0000; data[1442] = 16'h0000; data[1443] = 16'h0000; data[1444] = 16'h0000; data[1445] = 16'h0000; data[1446] = 16'h0000; data[1447] =
16'h0000; data[1448] = 16'h574b; data[1449] = 16'h52dc; data[1450] = 16'h460d; data[1451] = 16'h5249; data[1452] = 16'h55f4; data[1453] = 16'h4f70; data[1454] = 16'h0000; data[1455] = 16'h5416; data[1456] = 16'h5861; data[1457] = 16'h50ea; data[1458] = 16'h4d19; data[1459] = 16'h50a8; data[1460] = 16'h5579; data[1461] = 16'h4dc1; data[1462] = 16'h52d9; data[1463] = 16'h56b5; data[1464] = 16'h0000; data[1465] = 16'h0000; data[1466] = 16'h0000; data[1467] = 16'h0000; data[1468] = 16'h0000; data[1469]
= 16'h0000; data[1470] = 16'h0000; data[1471] = 16'h0000; data[1472] = 16'h5933; data[1473] = 16'h51fb; data[1474] = 16'h5266; data[1475] = 16'h522f; data[1476] = 16'h56d9; data[1477] = 16'h4d6e; data[1478] = 16'h0000; data[1479] = 16'h54be; data[1480] = 16'h58f1; data[1481] = 16'h52f5;
data[1482] = 16'h5718; data[1483] = 16'h5331; data[1484] = 16'h566d; data[1485] = 16'h4d47; data[1486] = 16'h4ff9; data[1487] = 16'h560c; data[1488] = 16'h0000; data[1489] = 16'h0000; data[1490] = 16'h0000; data[1491] = 16'h0000; data[1492] = 16'h0000; data[1493] = 16'h0000; data[1494] = 16'h0000; data[1495] = 16'h0000; data[1496] = 16'h56a5; data[1497] = 16'h5597; data[1498] = 16'h56e2; data[1499] = 16'h5155; data[1500] = 16'h56b8; data[1501] = 16'h4d9e; data[1502] = 16'h5786; data[1503] = 16'h4ff1; data[1504] = 16'h5440; data[1505] = 16'h58ea; data[1506] = 16'h58be; data[1507] = 16'h534f; data[1508] = 16'h561b; data[1509] = 16'h4bb1; data[1510] = 16'h58a9; data[1511] = 16'h0000; data[1512] = 16'h0000; data[1513] = 16'h0000; data[1514] = 16'h0000; data[1515] = 16'h0000; data[1516] = 16'h0000; data[1517] = 16'h0000; data[1518] = 16'h0000; data[1519] =
16'h0000; data[1520] = 16'h5457; data[1521] = 16'h5582; data[1522] = 16'h56d3; data[1523] = 16'h534b; data[1524] = 16'h568f; data[1525] = 16'h4940; data[1526] = 16'h544c; data[1527] = 16'h35c0; data[1528] = 16'h5029; data[1529] = 16'h59be; data[1530] = 16'h0000; data[1531] = 16'h5090; data[1532] = 16'h5722; data[1533] = 16'h0000; data[1534] = 16'h5690; data[1535] = 16'h5069; data[1536] = 16'h0000; data[1537] = 16'h0000; data[1538] = 16'h0000; data[1539] = 16'h0000; data[1540] = 16'h0000; data[1541]
= 16'h0000; data[1542] = 16'h0000; data[1543] = 16'h0000; data[1544] = 16'h5790; data[1545] = 16'h529d; data[1546] = 16'h4c5a; data[1547] = 16'h4fc3; data[1548] = 16'h5590; data[1549] = 16'h4d8b; data[1550] = 16'h427e; data[1551] = 16'h5602; data[1552] = 16'h4e4a; data[1553] = 16'h5626;
data[1554] = 16'h0000; data[1555] = 16'h49d2; data[1556] = 16'h5792; data[1557] = 16'h3e64; data[1558] = 16'h546c; data[1559] = 16'h57d8; data[1560] = 16'h0000; data[1561] = 16'h0000; data[1562] = 16'h0000; data[1563] = 16'h0000; data[1564] = 16'h0000; data[1565] = 16'h0000; data[1566] = 16'h0000; data[1567] = 16'h0000; data[1568] = 16'h5450; data[1569] = 16'h0000; data[1570] = 16'h54fb; data[1571] = 16'h493b; data[1572] = 16'h542b; data[1573] = 16'h4b07; data[1574] = 16'h0000; data[1575] = 16'h555d; data[1576] = 16'h4cc7; data[1577] = 16'h0000; data[1578] = 16'h55b9; data[1579] = 16'h4958; data[1580] = 16'h54cd; data[1581] = 16'h48e3; data[1582] = 16'h51a6; data[1583] = 16'h54b6; data[1584] = 16'h0000; data[1585] = 16'h0000; data[1586] = 16'h0000; data[1587] = 16'h0000; data[1588] = 16'h0000; data[1589] = 16'h0000; data[1590] = 16'h0000; data[1591] =
16'h0000; data[1592] = 16'h5362; data[1593] = 16'h5390; data[1594] = 16'h5849; data[1595] = 16'h4d32; data[1596] = 16'h5848; data[1597] = 16'h48bc; data[1598] = 16'h0000; data[1599] = 16'h52d5; data[1600] = 16'h5373; data[1601] = 16'h5068; data[1602] = 16'h5551; data[1603] = 16'h4a04; data[1604] = 16'h5818; data[1605] = 16'h4a68; data[1606] = 16'h526a; data[1607] = 16'h5400; data[1608] = 16'h0000; data[1609] = 16'h0000; data[1610] = 16'h0000; data[1611] = 16'h0000; data[1612] = 16'h0000; data[1613]
= 16'h0000; data[1614] = 16'h0000; data[1615] = 16'h0000; data[1616] = 16'h5535; data[1617] = 16'h53f5; data[1618] = 16'h5060; data[1619] = 16'h4d10; data[1620] = 16'h5818; data[1621] = 16'h4f0c; data[1622] = 16'h4bde; data[1623] = 16'h4a7f; data[1624] = 16'h5533; data[1625] = 16'h53d3;
data[1626] = 16'h5472; data[1627] = 16'h4cdb; data[1628] = 16'h577c; data[1629] = 16'h4d04; data[1630] = 16'h54c7; data[1631] = 16'h4be2; data[1632] = 16'h0000; data[1633] = 16'h0000; data[1634] = 16'h0000; data[1635] = 16'h0000; data[1636] = 16'h0000; data[1637] = 16'h0000; data[1638] = 16'h0000; data[1639] = 16'h0000; data[1640] = 16'h5517; data[1641] = 16'h5662; data[1642] = 16'h0000; data[1643] = 16'h525c; data[1644] = 16'h57c6; data[1645] = 16'h52cc; data[1646] = 16'h5516; data[1647] = 16'h53da; data[1648] = 16'h54e1; data[1649] = 16'h553c; data[1650] = 16'h4ff3; data[1651] = 16'h4ea2; data[1652] = 16'h5707; data[1653] = 16'h4f99; data[1654] = 16'h4e86; data[1655] = 16'h4f80; data[1656] = 16'h0000; data[1657] = 16'h0000; data[1658] = 16'h0000; data[1659] = 16'h0000; data[1660] = 16'h0000; data[1661] = 16'h0000; data[1662] = 16'h0000; data[1663] =
16'h0000; data[1664] = 16'h565a; data[1665] = 16'h5468; data[1666] = 16'h4cd5; data[1667] = 16'h547d; data[1668] = 16'h5750; data[1669] = 16'h4ed8; data[1670] = 16'h519c; data[1671] = 16'h54c7; data[1672] = 16'h55e2; data[1673] = 16'h5446; data[1674] = 16'h0000; data[1675] = 16'h509e; data[1676] = 16'h56fd; data[1677] = 16'h4d47; data[1678] = 16'h4c54; data[1679] = 16'h5759; data[1680] = 16'h0000; data[1681] = 16'h0000; data[1682] = 16'h0000; data[1683] = 16'h0000; data[1684] = 16'h0000; data[1685]
= 16'h0000; data[1686] = 16'h0000; data[1687] = 16'h0000; data[1688] = 16'h5830; data[1689] = 16'h5488; data[1690] = 16'h568e; data[1691] = 16'h5499; data[1692] = 16'h5804; data[1693] = 16'h4e52; data[1694] = 16'h0000; data[1695] = 16'h534d; data[1696] = 16'h5574; data[1697] = 16'h0000;
data[1698] = 16'h4f07; data[1699] = 16'h504c; data[1700] = 16'h5788; data[1701] = 16'h5092; data[1702] = 16'h4f8f; data[1703] = 16'h57b2; data[1704] = 16'h0000; data[1705] = 16'h0000; data[1706] = 16'h0000; data[1707] = 16'h0000; data[1708] = 16'h0000; data[1709] = 16'h0000; data[1710] = 16'h0000; data[1711] = 16'h0000; data[1712] = 16'h575b; data[1713] = 16'h5471; data[1714] = 16'h51e3; data[1715] = 16'h4c24; data[1716] = 16'h58ac; data[1717] = 16'h4d66; data[1718] = 16'h0000; data[1719] = 16'h5680; data[1720] = 16'h527d; data[1721] = 16'h0000; data[1722] = 16'h5452; data[1723] = 16'h4f3f; data[1724] = 16'h58a9; data[1725] = 16'h4d2e; data[1726] = 16'h3984; data[1727] = 16'h55b1; data[1728] = 16'h0000; data[1729] = 16'h0000; data[1730] = 16'h0000; data[1731] = 16'h0000; data[1732] = 16'h0000; data[1733] = 16'h0000; data[1734] = 16'h0000; data[1735] =
16'h0000; data[1736] = 16'h54ff; data[1737] = 16'h43bb; data[1738] = 16'h5454; data[1739] = 16'h4fc9; data[1740] = 16'h589d; data[1741] = 16'h505a; data[1742] = 16'h0000; data[1743] = 16'h550e; data[1744] = 16'h51fb; data[1745] = 16'h43e3; data[1746] = 16'h523d; data[1747] = 16'h50ce; data[1748] = 16'h57f3; data[1749] = 16'h50d8; data[1750] = 16'h4d74; data[1751] = 16'h55b9; data[1752] = 16'h0000; data[1753] = 16'h0000; data[1754] = 16'h0000; data[1755] = 16'h0000; data[1756] = 16'h0000; data[1757]
= 16'h0000; data[1758] = 16'h0000; data[1759] = 16'h0000; data[1760] = 16'h5578; data[1761] = 16'h4bed; data[1762] = 16'h55d7; data[1763] = 16'h528a; data[1764] = 16'h5808; data[1765] = 16'h518f; data[1766] = 16'h0000; data[1767] = 16'h52e2; data[1768] = 16'h5410; data[1769] = 16'h497a;
data[1770] = 16'h52f9; data[1771] = 16'h50d5; data[1772] = 16'h5793; data[1773] = 16'h5089; data[1774] = 16'h486e; data[1775] = 16'h54fd; data[1776] = 16'h0000; data[1777] = 16'h0000; data[1778] = 16'h0000; data[1779] = 16'h0000; data[1780] = 16'h0000; data[1781] = 16'h0000; data[1782] = 16'h0000; data[1783] = 16'h0000; data[1784] = 16'h5299; data[1785] = 16'h4d36; data[1786] = 16'h52ef; data[1787] = 16'h5472; data[1788] = 16'h5808; data[1789] = 16'h4f52; data[1790] = 16'h4f5a; data[1791] = 16'h52fa; data[1792] = 16'h5237; data[1793] = 16'h54fe; data[1794] = 16'h5417; data[1795] = 16'h4eba; data[1796] = 16'h5884; data[1797] = 16'h4e11; data[1798] = 16'h5426; data[1799] = 16'h50e1; data[1800] = 16'h0000; data[1801] = 16'h0000; data[1802] = 16'h0000; data[1803] = 16'h0000; data[1804] = 16'h0000; data[1805] = 16'h0000; data[1806] = 16'h0000; data[1807] =
16'h0000; data[1808] = 16'h5178; data[1809] = 16'h4a81; data[1810] = 16'h521b; data[1811] = 16'h51c9; data[1812] = 16'h5878; data[1813] = 16'h4ffa; data[1814] = 16'h5413; data[1815] = 16'h5661; data[1816] = 16'h4df4; data[1817] = 16'h5821; data[1818] = 16'h531e; data[1819] = 16'h50e7; data[1820] = 16'h5863; data[1821] = 16'h4ff0; data[1822] = 16'h57f5; data[1823] = 16'h5318; data[1824] = 16'h0000; data[1825] = 16'h0000; data[1826] = 16'h0000; data[1827] = 16'h0000; data[1828] = 16'h0000; data[1829]
= 16'h0000; data[1830] = 16'h0000; data[1831] = 16'h0000; data[1832] = 16'h559a; data[1833] = 16'h4902; data[1834] = 16'h5524; data[1835] = 16'h51d3; data[1836] = 16'h584a; data[1837] = 16'h521e; data[1838] = 16'h5296; data[1839] = 16'h57b2; data[1840] = 16'h5375; data[1841] = 16'h569e;
data[1842] = 16'h5961; data[1843] = 16'h55b3; data[1844] = 16'h5963; data[1845] = 16'h4f0a; data[1846] = 16'h577b; data[1847] = 16'h53e2; data[1848] = 16'h0000; data[1849] = 16'h0000; data[1850] = 16'h0000; data[1851] = 16'h0000; data[1852] = 16'h0000; data[1853] = 16'h0000; data[1854] = 16'h0000; data[1855] = 16'h0000; data[1856] = 16'h56cd; data[1857] = 16'h4612; data[1858] = 16'h5923; data[1859] = 16'h51ce; data[1860] = 16'h585b; data[1861] = 16'h5268; data[1862] = 16'h4f4a; data[1863] = 16'h54eb; data[1864] = 16'h5664; data[1865] = 16'h535e; data[1866] = 16'h5660; data[1867] = 16'h561e; data[1868] = 16'h58d9; data[1869] = 16'h4f89; data[1870] = 16'h55cb; data[1871] = 16'h55a7; data[1872] = 16'h0000; data[1873] = 16'h0000; data[1874] = 16'h0000; data[1875] = 16'h0000; data[1876] = 16'h0000; data[1877] = 16'h0000; data[1878] = 16'h0000; data[1879] =
16'h0000; data[1880] = 16'h55f5; data[1881] = 16'h50ef; data[1882] = 16'h583f; data[1883] = 16'h4d0e; data[1884] = 16'h582d; data[1885] = 16'h4ec6; data[1886] = 16'h4e9a; data[1887] = 16'h4d7e; data[1888] = 16'h568e; data[1889] = 16'h4f0f; data[1890] = 16'h585f; data[1891] = 16'h5256; data[1892] = 16'h5831; data[1893] = 16'h4d89; data[1894] = 16'h529d; data[1895] = 16'h5196; data[1896] = 16'h0000; data[1897] = 16'h0000; data[1898] = 16'h0000; data[1899] = 16'h0000; data[1900] = 16'h0000; data[1901]
= 16'h0000; data[1902] = 16'h0000; data[1903] = 16'h0000; data[1904] = 16'h5596; data[1905] = 16'h5379; data[1906] = 16'h55c2; data[1907] = 16'h4f14; data[1908] = 16'h56fa; data[1909] = 16'h50b7; data[1910] = 16'h4f2e; data[1911] = 16'h48d2; data[1912] = 16'h5554; data[1913] = 16'h53cf;
data[1914] = 16'h51a2; data[1915] = 16'h521f; data[1916] = 16'h574d; data[1917] = 16'h4fbc; data[1918] = 16'h0000; data[1919] = 16'h51f1; data[1920] = 16'h0000; data[1921] = 16'h0000; data[1922] = 16'h0000; data[1923] = 16'h0000; data[1924] = 16'h0000; data[1925] = 16'h0000; data[1926] = 16'h0000; data[1927] = 16'h0000; data[1928] = 16'h55ed; data[1929] = 16'h5500; data[1930] = 16'h54b8; data[1931] = 16'h4f08; data[1932] = 16'h56c8; data[1933] = 16'h4ebb; data[1934] = 16'h0000; data[1935] = 16'h4787; data[1936] = 16'h55d6; data[1937] = 16'h53a6; data[1938] = 16'h4e78; data[1939] = 16'h4ee8; data[1940] = 16'h56f8; data[1941] = 16'h4e50; data[1942] = 16'h0000; data[1943] = 16'h5157; data[1944] = 16'h0000; data[1945] = 16'h0000; data[1946] = 16'h0000; data[1947] = 16'h0000; data[1948] = 16'h0000; data[1949] = 16'h0000; data[1950] = 16'h0000; data[1951] =
16'h0000; data[1952] = 16'h5633; data[1953] = 16'h5679; data[1954] = 16'h0000; data[1955] = 16'h4e58; data[1956] = 16'h5820; data[1957] = 16'h4db0; data[1958] = 16'h5032; data[1959] = 16'h536d; data[1960] = 16'h5605; data[1961] = 16'h522b; data[1962] = 16'h45e1; data[1963] = 16'h4a9c; data[1964] = 16'h570c; data[1965] = 16'h4ec2; data[1966] = 16'h0000; data[1967] = 16'h525f; data[1968] = 16'h0000; data[1969] = 16'h0000; data[1970] = 16'h0000; data[1971] = 16'h0000; data[1972] = 16'h0000; data[1973]
= 16'h0000; data[1974] = 16'h0000; data[1975] = 16'h0000; data[1976] = 16'h54f8; data[1977] = 16'h502f; data[1978] = 16'h0000; data[1979] = 16'h4cc6; data[1980] = 16'h57f7; data[1981] = 16'h4e9a; data[1982] = 16'h52f0; data[1983] = 16'h5560; data[1984] = 16'h55b7; data[1985] = 16'h506a;
data[1986] = 16'h5149; data[1987] = 16'h4e49; data[1988] = 16'h566a; data[1989] = 16'h4fae; data[1990] = 16'h5214; data[1991] = 16'h5322; data[1992] = 16'h0000; data[1993] = 16'h0000; data[1994] = 16'h0000; data[1995] = 16'h0000; data[1996] = 16'h0000; data[1997] = 16'h0000; data[1998] = 16'h0000; data[1999] = 16'h0000; data[2000] = 16'h525b; data[2001] = 16'h4c1c; data[2002] = 16'h55b5; data[2003] = 16'h4bcf; data[2004] = 16'h578e; data[2005] = 16'h508d; data[2006] = 16'h528b; data[2007] = 16'h512c; data[2008] = 16'h55fb; data[2009] = 16'h4f8a; data[2010] = 16'h54b2; data[2011] = 16'h5091; data[2012] = 16'h5769; data[2013] = 16'h4e87; data[2014] = 16'h514f; data[2015] = 16'h5131; data[2016] = 16'h0000; data[2017] = 16'h0000; data[2018] = 16'h0000; data[2019] = 16'h0000; data[2020] = 16'h0000; data[2021] = 16'h0000; data[2022] = 16'h0000; data[2023] =
16'h0000; data[2024] = 16'h54ee; data[2025] = 16'h4c3a; data[2026] = 16'h5006; data[2027] = 16'h4a05; data[2028] = 16'h5804; data[2029] = 16'h5127; data[2030] = 16'h4fae; data[2031] = 16'h58e6; data[2032] = 16'h5534; data[2033] = 16'h4518; data[2034] = 16'h5546; data[2035] = 16'h4939; data[2036] = 16'h584e; data[2037] = 16'h502e; data[2038] = 16'h4d8b; data[2039] = 16'h5882; data[2040] = 16'h0000; data[2041] = 16'h0000; data[2042] = 16'h0000; data[2043] = 16'h0000; data[2044] = 16'h0000; data[2045]
= 16'h0000; data[2046] = 16'h0000; data[2047] = 16'h0000; data[2048] = 16'h55b1; data[2049] = 16'h0000; data[2050] = 16'h56df; data[2051] = 16'h486f; data[2052] = 16'h57b0; data[2053] = 16'h4cb8; data[2054] = 16'h4ede; data[2055] = 16'h56f6; data[2056] = 16'h54b0; data[2057] = 16'h46d7;
data[2058] = 16'h5871; data[2059] = 16'h4eac; data[2060] = 16'h5813; data[2061] = 16'h51f1; data[2062] = 16'h5298; data[2063] = 16'h5734; data[2064] = 16'h0000; data[2065] = 16'h0000; data[2066] = 16'h0000; data[2067] = 16'h0000; data[2068] = 16'h0000; data[2069] = 16'h0000; data[2070] = 16'h0000; data[2071] = 16'h0000; data[2072] = 16'h540e; data[2073] = 16'h4438; data[2074] = 16'h51c0; data[2075] = 16'h4b16; data[2076] = 16'h567e; data[2077] = 16'h4dec; data[2078] = 16'h0000; data[2079] = 16'h55ef; data[2080] = 16'h5ab4; data[2081] = 16'h4da2; data[2082] = 16'h0000; data[2083] = 16'h506b; data[2084] = 16'h564a; data[2085] = 16'h54db; data[2086] = 16'h0000; data[2087] = 16'h5b32; data[2088] = 16'h0000; data[2089] = 16'h0000; data[2090] = 16'h0000; data[2091] = 16'h0000; data[2092] = 16'h0000; data[2093] = 16'h0000; data[2094] = 16'h0000; data[2095] =
16'h0000; data[2096] = 16'h59b1; data[2097] = 16'h424f; data[2098] = 16'h4caa; data[2099] = 16'h4cfc; data[2100] = 16'h560c; data[2101] = 16'h51f6; data[2102] = 16'h0000; data[2103] = 16'h566b; data[2104] = 16'h5c5f; data[2105] = 16'h4f1c; data[2106] = 16'h55b3; data[2107] = 16'h538c; data[2108] = 16'h5728; data[2109] = 16'h546f; data[2110] = 16'h0000; data[2111] = 16'h5edd; data[2112] = 16'h0000; data[2113] = 16'h0000; data[2114] = 16'h0000; data[2115] = 16'h0000; data[2116] = 16'h0000; data[2117]
= 16'h0000; data[2118] = 16'h0000; data[2119] = 16'h0000; data[2120] = 16'h5c9e; data[2121] = 16'h4d10; data[2122] = 16'h51ee; data[2123] = 16'h5372; data[2124] = 16'h56e1; data[2125] = 16'h5434; data[2126] = 16'h0000; data[2127] = 16'h5e1d; data[2128] = 16'h5c9b; data[2129] = 16'h4f9e;
data[2130] = 16'h559b; data[2131] = 16'h5315; data[2132] = 16'h5578; data[2133] = 16'h554e; data[2134] = 16'h0000; data[2135] = 16'h5f27; data[2136] = 16'h0000; data[2137] = 16'h0000; data[2138] = 16'h0000; data[2139] = 16'h0000; data[2140] = 16'h0000; data[2141] = 16'h0000; data[2142] = 16'h0000; data[2143] = 16'h0000; data[2144] = 16'h5c98; data[2145] = 16'h4cc4; data[2146] = 16'h56ee; data[2147] = 16'h541e; data[2148] = 16'h5672; data[2149] = 16'h5333; data[2150] = 16'h0000; data[2151] = 16'h5ef8; data[2152] = 16'h5899; data[2153] = 16'h4ce4; data[2154] = 16'h5837; data[2155] = 16'h4ccb; data[2156] = 16'h5090; data[2157] = 16'h5469; data[2158] = 16'h0000; data[2159] = 16'h5f1e; data[2160] = 16'h0000; data[2161] = 16'h0000; data[2162] = 16'h0000; data[2163] = 16'h0000; data[2164] = 16'h0000; data[2165] = 16'h0000; data[2166] = 16'h0000; data[2167] =
16'h0000; data[2168] = 16'h5d77; data[2169] = 16'h0000; data[2170] = 16'h5cf4; data[2171] = 16'h55d1; data[2172] = 16'h58a4; data[2173] = 16'h50f5; data[2174] = 16'h0000; data[2175] = 16'h5d11; data[2176] = 16'h55b4; data[2177] = 16'h40f2; data[2178] = 16'h5bc0; data[2179] = 16'h526e; data[2180] = 16'h5371; data[2181] = 16'h4d60; data[2182] = 16'h0000; data[2183] = 16'h5dc3; data[2184] = 16'h0000; data[2185] = 16'h0000; data[2186] = 16'h0000; data[2187] = 16'h0000; data[2188] = 16'h0000; data[2189]
= 16'h0000; data[2190] = 16'h0000; data[2191] = 16'h0000; data[2192] = 16'h5c64; data[2193] = 16'h0000; data[2194] = 16'h5cb0; data[2195] = 16'h5816; data[2196] = 16'h5965; data[2197] = 16'h5263; data[2198] = 16'h0000; data[2199] = 16'h5c58; data[2200] = 16'h5c6e; data[2201] = 16'h0000;
data[2202] = 16'h5cf8; data[2203] = 16'h54d8; data[2204] = 16'h55a2; data[2205] = 16'h4f24; data[2206] = 16'h0000; data[2207] = 16'h5cf9; data[2208] = 16'h0000; data[2209] = 16'h0000; data[2210] = 16'h0000; data[2211] = 16'h0000; data[2212] = 16'h0000; data[2213] = 16'h0000; data[2214] = 16'h0000; data[2215] = 16'h0000; data[2216] = 16'h5bca; data[2217] = 16'h0000; data[2218] = 16'h5931; data[2219] = 16'h54ef; data[2220] = 16'h57c1; data[2221] = 16'h518e; data[2222] = 16'h0000; data[2223] = 16'h587c; data[2224] = 16'h5c90; data[2225] = 16'h0000; data[2226] = 16'h5db5; data[2227] = 16'h5898; data[2228] = 16'h567d; data[2229] = 16'h4eb0; data[2230] = 16'h0000; data[2231] = 16'h5c7c; data[2232] = 16'h0000; data[2233] = 16'h0000; data[2234] = 16'h0000; data[2235] = 16'h0000; data[2236] = 16'h0000; data[2237] = 16'h0000; data[2238] = 16'h0000; data[2239] =
16'h0000; data[2240] = 16'h5639; data[2241] = 16'h0000; data[2242] = 16'h5847; data[2243] = 16'h5630; data[2244] = 16'h5796; data[2245] = 16'h4e08; data[2246] = 16'h4560; data[2247] = 16'h582d; data[2248] = 16'h5af8; data[2249] = 16'h0000; data[2250] = 16'h5d2e; data[2251] = 16'h5898; data[2252] = 16'h5906; data[2253] = 16'h4bed; data[2254] = 16'h0000; data[2255] = 16'h5c4b; data[2256] = 16'h0000; data[2257] = 16'h0000; data[2258] = 16'h0000; data[2259] = 16'h0000; data[2260] = 16'h0000; data[2261]
= 16'h0000; data[2262] = 16'h0000; data[2263] = 16'h0000; data[2264] = 16'h5379; data[2265] = 16'h0000; data[2266] = 16'h572b; data[2267] = 16'h5019; data[2268] = 16'h572e; data[2269] = 16'h4dea; data[2270] = 16'h4311; data[2271] = 16'h5853; data[2272] = 16'h5410; data[2273] = 16'h0000;
data[2274] = 16'h5881; data[2275] = 16'h5406; data[2276] = 16'h587c; data[2277] = 16'h4df2; data[2278] = 16'h0000; data[2279] = 16'h58a5; data[2280] = 16'h0000; data[2281] = 16'h0000; data[2282] = 16'h0000; data[2283] = 16'h0000; data[2284] = 16'h0000; data[2285] = 16'h0000; data[2286] = 16'h0000; data[2287] = 16'h0000; data[2288] = 16'h50e5; data[2289] = 16'h0000; data[2290] = 16'h5632; data[2291] = 16'h500a; data[2292] = 16'h576d; data[2293] = 16'h4e3a; data[2294] = 16'h0000; data[2295] = 16'h5646; data[2296] = 16'h5321; data[2297] = 16'h0000; data[2298] = 16'h582a; data[2299] = 16'h50a3; data[2300] = 16'h5783; data[2301] = 16'h4d4c; data[2302] = 16'h4442; data[2303] = 16'h5680; data[2304] = 16'h0000; data[2305] = 16'h0000; data[2306] = 16'h0000; data[2307] = 16'h0000; data[2308] = 16'h0000; data[2309] = 16'h0000; data[2310] = 16'h0000; data[2311] =
16'h0000; data[2312] = 16'h5212; data[2313] = 16'h0000; data[2314] = 16'h556e; data[2315] = 16'h4f4b; data[2316] = 16'h5753; data[2317] = 16'h4c99; data[2318] = 16'h4098; data[2319] = 16'h583e; data[2320] = 16'h51c9; data[2321] = 16'h399a; data[2322] = 16'h5438; data[2323] = 16'h4ec0; data[2324] = 16'h56f9; data[2325] = 16'h4df0; data[2326] = 16'h4444; data[2327] = 16'h5836; data[2328] = 16'h0000; data[2329] = 16'h0000; data[2330] = 16'h0000; data[2331] = 16'h0000; data[2332] = 16'h0000; data[2333]
= 16'h0000; data[2334] = 16'h0000; data[2335] = 16'h0000; data[2336] = 16'h51df; data[2337] = 16'h0000; data[2338] = 16'h5808; data[2339] = 16'h5088; data[2340] = 16'h5806; data[2341] = 16'h4d09; data[2342] = 16'h4295; data[2343] = 16'h56f8; data[2344] = 16'h512e; data[2345] = 16'h3a10;
data[2346] = 16'h5685; data[2347] = 16'h4fbc; data[2348] = 16'h574b; data[2349] = 16'h4eda; data[2350] = 16'h4b48; data[2351] = 16'h566a; data[2352] = 16'h0000; data[2353] = 16'h0000; data[2354] = 16'h0000; data[2355] = 16'h0000; data[2356] = 16'h0000; data[2357] = 16'h0000; data[2358] = 16'h0000; data[2359] = 16'h0000; data[2360] = 16'h5044; data[2361] = 16'h3ecc; data[2362] = 16'h54cd; data[2363] = 16'h4f09; data[2364] = 16'h57a1; data[2365] = 16'h4e99; data[2366] = 16'h4f80; data[2367] = 16'h5340; data[2368] = 16'h53f1; data[2369] = 16'h41cf; data[2370] = 16'h5421; data[2371] = 16'h4e32; data[2372] = 16'h57e0; data[2373] = 16'h4f49; data[2374] = 16'h0000; data[2375] = 16'h5596; data[2376] = 16'h0000; data[2377] = 16'h0000; data[2378] = 16'h0000; data[2379] = 16'h0000; data[2380] = 16'h0000; data[2381] = 16'h0000; data[2382] = 16'h0000; data[2383] =
16'h0000; data[2384] = 16'h5367; data[2385] = 16'h46c4; data[2386] = 16'h4d7f; data[2387] = 16'h4f33; data[2388] = 16'h5701; data[2389] = 16'h4e57; data[2390] = 16'h4816; data[2391] = 16'h55d1; data[2392] = 16'h5179; data[2393] = 16'h45a1; data[2394] = 16'h53b2; data[2395] = 16'h4ae1; data[2396] = 16'h5702; data[2397] = 16'h4f49; data[2398] = 16'h0000; data[2399] = 16'h55a2; data[2400] = 16'h0000; data[2401] = 16'h0000; data[2402] = 16'h0000; data[2403] = 16'h0000; data[2404] = 16'h0000; data[2405]
= 16'h0000; data[2406] = 16'h0000; data[2407] = 16'h0000; data[2408] = 16'h54ba; data[2409] = 16'h44c7; data[2410] = 16'h521d; data[2411] = 16'h4e5e; data[2412] = 16'h5764; data[2413] = 16'h4e28; data[2414] = 16'h0000; data[2415] = 16'h57f9; data[2416] = 16'h4d38; data[2417] = 16'h4358;
data[2418] = 16'h52cd; data[2419] = 16'h49f2; data[2420] = 16'h56e8; data[2421] = 16'h4e08; data[2422] = 16'h5079; data[2423] = 16'h57c0; data[2424] = 16'h0000; data[2425] = 16'h0000; data[2426] = 16'h0000; data[2427] = 16'h0000; data[2428] = 16'h0000; data[2429] = 16'h0000; data[2430] = 16'h0000; data[2431] = 16'h0000; data[2432] = 16'h5431; data[2433] = 16'h0000; data[2434] = 16'h55f2; data[2435] = 16'h4558; data[2436] = 16'h57ac; data[2437] = 16'h4df2; data[2438] = 16'h4aa8; data[2439] = 16'h57cd; data[2440] = 16'h4ca8; data[2441] = 16'h4040; data[2442] = 16'h5555; data[2443] = 16'h4dd8; data[2444] = 16'h578b; data[2445] = 16'h4e3b; data[2446] = 16'h52be; data[2447] = 16'h56cb; data[2448] = 16'h0000; data[2449] = 16'h0000; data[2450] = 16'h0000; data[2451] = 16'h0000; data[2452] = 16'h0000; data[2453] = 16'h0000; data[2454] = 16'h0000; data[2455] =
16'h0000; data[2456] = 16'h50d2; data[2457] = 16'h0000; data[2458] = 16'h551d; data[2459] = 16'h45cc; data[2460] = 16'h5766; data[2461] = 16'h4f7d; data[2462] = 16'h4216; data[2463] = 16'h5555; data[2464] = 16'h5097; data[2465] = 16'h4182; data[2466] = 16'h53eb; data[2467] = 16'h4d96; data[2468] = 16'h56c0; data[2469] = 16'h5040; data[2470] = 16'h49a0; data[2471] = 16'h550c; data[2472] = 16'h0000; data[2473] = 16'h0000; data[2474] = 16'h0000; data[2475] = 16'h0000; data[2476] = 16'h0000; data[2477]
= 16'h0000; data[2478] = 16'h0000; data[2479] = 16'h0000; data[2480] = 16'h5312; data[2481] = 16'h4937; data[2482] = 16'h5036; data[2483] = 16'h4a7a; data[2484] = 16'h5732; data[2485] = 16'h5012; data[2486] = 16'h2ccc; data[2487] = 16'h5870; data[2488] = 16'h5176; data[2489] = 16'h4513;
data[2490] = 16'h53f3; data[2491] = 16'h4981; data[2492] = 16'h570b; data[2493] = 16'h4df7; data[2494] = 16'h4ca1; data[2495] = 16'h573d; data[2496] = 16'h0000; data[2497] = 16'h0000; data[2498] = 16'h0000; data[2499] = 16'h0000; data[2500] = 16'h0000; data[2501] = 16'h0000; data[2502] = 16'h0000; data[2503] = 16'h0000; data[2504] = 16'h5371; data[2505] = 16'h0000; data[2506] = 16'h55d1; data[2507] = 16'h4b14; data[2508] = 16'h5771; data[2509] = 16'h4e66; data[2510] = 16'h480a; data[2511] = 16'h586b; data[2512] = 16'h505c; data[2513] = 16'h0000; data[2514] = 16'h5727; data[2515] = 16'h4d9c; data[2516] = 16'h56f5; data[2517] = 16'h4d93; data[2518] = 16'h4edd; data[2519] = 16'h569e; data[2520] = 16'h0000; data[2521] = 16'h0000; data[2522] = 16'h0000; data[2523] = 16'h0000; data[2524] = 16'h0000; data[2525] = 16'h0000; data[2526] = 16'h0000; data[2527] =
16'h0000; data[2528] = 16'h4df1; data[2529] = 16'h4886; data[2530] = 16'h580a; data[2531] = 16'h4ca3; data[2532] = 16'h5833; data[2533] = 16'h501c; data[2534] = 16'h501a; data[2535] = 16'h556e; data[2536] = 16'h5377; data[2537] = 16'h4702; data[2538] = 16'h5549; data[2539] = 16'h4ae6; data[2540] = 16'h585a; data[2541] = 16'h4f35; data[2542] = 16'h0000; data[2543] = 16'h54bc; data[2544] = 16'h0000; data[2545] = 16'h0000; data[2546] = 16'h0000; data[2547] = 16'h0000; data[2548] = 16'h0000; data[2549]
= 16'h0000; data[2550] = 16'h0000; data[2551] = 16'h0000; data[2552] = 16'h4cbc; data[2553] = 16'h4d16; data[2554] = 16'h5195; data[2555] = 16'h496d; data[2556] = 16'h57ac; data[2557] = 16'h504f; data[2558] = 16'h5271; data[2559] = 16'h56f1; data[2560] = 16'h5400; data[2561] = 16'h4a97;
data[2562] = 16'h529a; data[2563] = 16'h45da; data[2564] = 16'h580b; data[2565] = 16'h511d; data[2566] = 16'h0000; data[2567] = 16'h55f3; data[2568] = 16'h0000; data[2569] = 16'h0000; data[2570] = 16'h0000; data[2571] = 16'h0000; data[2572] = 16'h0000; data[2573] = 16'h0000; data[2574] = 16'h0000; data[2575] = 16'h0000; data[2576] = 16'h4a11; data[2577] = 16'h3a5c; data[2578] = 16'h54f0; data[2579] = 16'h49e1; data[2580] = 16'h56d1; data[2581] = 16'h4ef8; data[2582] = 16'h5495; data[2583] = 16'h5759; data[2584] = 16'h5150; data[2585] = 16'h459c; data[2586] = 16'h526b; data[2587] = 16'h4c23; data[2588] = 16'h56a6; data[2589] = 16'h4fac; data[2590] = 16'h4e85; data[2591] = 16'h5418; data[2592] = 16'h0000; data[2593] = 16'h0000; data[2594] = 16'h0000; data[2595] = 16'h0000; data[2596] = 16'h0000; data[2597] = 16'h0000; data[2598] = 16'h0000; data[2599] =
16'h0000; data[2600] = 16'h5200; data[2601] = 16'h0000; data[2602] = 16'h5624; data[2603] = 16'h48a7; data[2604] = 16'h5869; data[2605] = 16'h4d1a; data[2606] = 16'h511a; data[2607] = 16'h5643; data[2608] = 16'h5211; data[2609] = 16'h49c3; data[2610] = 16'h5010; data[2611] = 16'h4a24; data[2612] = 16'h57b9; data[2613] = 16'h4d92; data[2614] = 16'h4bf1; data[2615] = 16'h5673; data[2616] = 16'h0000; data[2617] = 16'h0000; data[2618] = 16'h0000; data[2619] = 16'h0000; data[2620] = 16'h0000; data[2621]
= 16'h0000; data[2622] = 16'h0000; data[2623] = 16'h0000; data[2624] = 16'h4f89; data[2625] = 16'h4718; data[2626] = 16'h5150; data[2627] = 16'h4a19; data[2628] = 16'h57ff; data[2629] = 16'h4ef1; data[2630] = 16'h508f; data[2631] = 16'h5805; data[2632] = 16'h4ef2; data[2633] = 16'h43ae;
data[2634] = 16'h531d; data[2635] = 16'h4a5e; data[2636] = 16'h57d1; data[2637] = 16'h501f; data[2638] = 16'h4c08; data[2639] = 16'h5697; data[2640] = 16'h0000; data[2641] = 16'h0000; data[2642] = 16'h0000; data[2643] = 16'h0000; data[2644] = 16'h0000; data[2645] = 16'h0000; data[2646] = 16'h0000; data[2647] = 16'h0000; data[2648] = 16'h50aa; data[2649] = 16'h4250; data[2650] = 16'h55c0; data[2651] = 16'h4aec; data[2652] = 16'h5799; data[2653] = 16'h4f90; data[2654] = 16'h4dc3; data[2655] = 16'h56df; data[2656] = 16'h50c6; data[2657] = 16'h4298; data[2658] = 16'h5572; data[2659] = 16'h4b15; data[2660] = 16'h575c; data[2661] = 16'h5040; data[2662] = 16'h4c9f; data[2663] = 16'h56c7; data[2664] = 16'h0000; data[2665] = 16'h0000; data[2666] = 16'h0000; data[2667] = 16'h0000; data[2668] = 16'h0000; data[2669] = 16'h0000; data[2670] = 16'h0000; data[2671] =
16'h0000; data[2672] = 16'h508d; data[2673] = 16'h4412; data[2674] = 16'h551c; data[2675] = 16'h4b48; data[2676] = 16'h5754; data[2677] = 16'h50af; data[2678] = 16'h51a3; data[2679] = 16'h5793; data[2680] = 16'h50c0; data[2681] = 16'h0000; data[2682] = 16'h555e; data[2683] = 16'h4d1e; data[2684] = 16'h56d4; data[2685] = 16'h4e66; data[2686] = 16'h4cb2; data[2687] = 16'h567f; data[2688] = 16'h0000; data[2689] = 16'h0000; data[2690] = 16'h0000; data[2691] = 16'h0000; data[2692] = 16'h0000; data[2693]
= 16'h0000; data[2694] = 16'h0000; data[2695] = 16'h0000; data[2696] = 16'h507f; data[2697] = 16'h0000; data[2698] = 16'h5603; data[2699] = 16'h4ba0; data[2700] = 16'h5747; data[2701] = 16'h5090; data[2702] = 16'h50a5; data[2703] = 16'h5944; data[2704] = 16'h4b85; data[2705] = 16'h3902;
data[2706] = 16'h5509; data[2707] = 16'h4b5d; data[2708] = 16'h5771; data[2709] = 16'h4f0a; data[2710] = 16'h5266; data[2711] = 16'h590e; data[2712] = 16'h0000; data[2713] = 16'h0000; data[2714] = 16'h0000; data[2715] = 16'h0000; data[2716] = 16'h0000; data[2717] = 16'h0000; data[2718] = 16'h0000; data[2719] = 16'h0000; data[2720] = 16'h5448; data[2721] = 16'h0000; data[2722] = 16'h5849; data[2723] = 16'h4b23; data[2724] = 16'h58eb; data[2725] = 16'h4e53; data[2726] = 16'h0000; data[2727] = 16'h5896; data[2728] = 16'h4eae; data[2729] = 16'h3dc4; data[2730] = 16'h56e4; data[2731] = 16'h4d3a; data[2732] = 16'h581c; data[2733] = 16'h4fb9; data[2734] = 16'h501e; data[2735] = 16'h589c; data[2736] = 16'h0000; data[2737] = 16'h0000; data[2738] = 16'h0000; data[2739] = 16'h0000; data[2740] = 16'h0000; data[2741] = 16'h0000; data[2742] = 16'h0000; data[2743] =
16'h0000; data[2744] = 16'h5229; data[2745] = 16'h48ee; data[2746] = 16'h547a; data[2747] = 16'h4763; data[2748] = 16'h588a; data[2749] = 16'h5161; data[2750] = 16'h0000; data[2751] = 16'h58d7; data[2752] = 16'h4eb5; data[2753] = 16'h4150; data[2754] = 16'h56ec; data[2755] = 16'h4cfd; data[2756] = 16'h5897; data[2757] = 16'h509c; data[2758] = 16'h4c7b; data[2759] = 16'h5809; data[2760] = 16'h0000; data[2761] = 16'h0000; data[2762] = 16'h0000; data[2763] = 16'h0000; data[2764] = 16'h0000; data[2765]
= 16'h0000; data[2766] = 16'h0000; data[2767] = 16'h0000; data[2768] = 16'h0000; data[2769] = 16'h0000; data[2770] = 16'h0000; data[2771] = 16'h0000; data[2772] = 16'h0000; data[2773] = 16'h0000; data[2774] = 16'h0000; data[2775] = 16'h0000; data[2776] = 16'h0000; data[2777] = 16'h0000;
data[2778] = 16'h0000; data[2779] = 16'h0000; data[2780] = 16'h0000; data[2781] = 16'h0000; data[2782] = 16'h0000; data[2783] = 16'h0000;

weight[0] = 16'ha9bf; weight[1] = 16'h2a01; weight[2] = 16'ha6ab; weight[3] = 16'hac65; weight[4] = 16'h28c1; weight[5] = 16'h262c; weight[6] =
16'h2e83; weight[7] = 16'h2634; weight[8] = 16'h29ec; weight[9] = 16'ha220; weight[10] = 16'hb1db; weight[11] = 16'h2216; weight[12] = 16'h8eac; weight[13] = 16'h2469; weight[14] = 16'h251b; weight[15] = 16'h25ec; weight[16] = 16'h22bf; weight[17] = 16'ha1e9; weight[18] = 16'haffb; weight[19] = 16'h2480; weight[20] = 16'h294a; weight[21] = 16'ha9f4; weight[22] = 16'h2dcf; weight[23] = 16'haa8f; weight[24] = 16'hac4b; weight[25]
= 16'h2e3e; weight[26] = 16'h95db; weight[27] = 16'hae22; weight[28] = 16'h2aac; weight[29] = 16'h2ced; weight[30] = 16'hadb5; weight[31] = 16'h24fa; weight[32] = 16'hae4f; weight[33] = 16'h28a9; weight[34] = 16'h96bc; weight[35] = 16'h9ae4; weight[36] = 16'hb384; weight[37] = 16'hadd3;
weight[38] = 16'hb4b7; weight[39] = 16'hb02e; weight[40] = 16'h068f; weight[41] = 16'h2a89; weight[42] = 16'h979e; weight[43] = 16'h2bb3; weight[44] = 16'h3023; weight[45] = 16'h2436; weight[46] = 16'ha895; weight[47] = 16'h20a5; weight[48] = 16'h9f0b; weight[49] = 16'h2547; weight[50] = 16'haeb4; weight[51] = 16'hb002; weight[52] = 16'h263f; weight[53] = 16'h2ad9; weight[54] = 16'h2c98; weight[55] = 16'h269d; weight[56] = 16'h1c27; weight[57] = 16'haa0c; weight[58] = 16'hb085; weight[59] = 16'ha6f6; weight[60] = 16'ha8f2; weight[61] = 16'h2d91; weight[62] = 16'h2b1f; weight[63] = 16'ha05e; weight[64] = 16'h08b1; weight[65] = 16'h1dde; weight[66] = 16'ha743; weight[67] = 16'h9af5; weight[68] = 16'h2c34; weight[69] = 16'h1e94; weight[70] = 16'h30a0; weight[71] = 16'ha820; weight[72] = 16'ha127; weight[73] = 16'h29c3; weight[74] = 16'h2dee; weight[75] =
16'h2286; weight[76] = 16'h2980; weight[77] = 16'haa78; weight[78] = 16'h244b; weight[79] = 16'h2902; weight[80] = 16'ha8f0; weight[81] = 16'ha8cc; weight[82] = 16'h1a01; weight[83] = 16'h2c25; weight[84] = 16'h13e1; weight[85] = 16'h2990; weight[86] = 16'ha68e; weight[87] = 16'h2850; weight[88] = 16'h2091; weight[89] = 16'h2e7d; weight[90] = 16'h28ca; weight[91] = 16'h2752; weight[92] = 16'h2e78; weight[93] = 16'ha9a9; weight[94] = 16'ha94d; weight[95] = 16'h2057; weight[96] = 16'hb0b0; weight[97]
= 16'ha4f7; weight[98] = 16'h2cae; weight[99] = 16'ha189; weight[100] =
16'ha9ae; weight[101] = 16'h28ae; weight[102] = 16'h219d; weight[103] =
16'h2f74; weight[104] = 16'hb7e8; weight[105] = 16'hb202; weight[106] =
16'h9bb6; weight[107] = 16'hb82a; weight[108] = 16'hb069; weight[109] =
16'ha9d7; weight[110] = 16'hb540; weight[111] = 16'haab9; weight[112] =
16'ha72a; weight[113] = 16'h2f4a; weight[114] = 16'h2139; weight[115] =
16'ha87f; weight[116] = 16'h2ee9; weight[117] = 16'h2d37; weight[118] =
16'hb0a1; weight[119] = 16'h2dc2; weight[120] = 16'h2367; weight[121] =
16'h2d90; weight[122] = 16'h28c0; weight[123] = 16'h308d; weight[124] =
16'h251e; weight[125] = 16'ha605; weight[126] = 16'h2c1d; weight[127] =
16'h2bda; weight[128] = 16'h2870; weight[129] = 16'h2419; weight[130] =
16'ha89b; weight[131] = 16'h3173; weight[132] = 16'ha1c0; weight[133] =
16'h1f98; weight[134] = 16'ha23d; weight[135] = 16'hace3; weight[136] =
16'h2b8f; weight[137] = 16'h323b; weight[138] = 16'h2b7e; weight[139] =
16'h3088; weight[140] = 16'h2e80; weight[141] = 16'h9b33; weight[142] =
16'h249c; weight[143] = 16'h295b; weight[144] = 16'hb004; weight[145] =
16'ha479; weight[146] = 16'h22c8; weight[147] = 16'h9195; weight[148] =
16'h2708; weight[149] = 16'h2dfe; weight[150] = 16'h2a61; weight[151] =
16'hac9f; weight[152] = 16'haf18; weight[153] = 16'h26ed; weight[154] =
16'hac97; weight[155] = 16'h28fd; weight[156] = 16'hae20; weight[157] =
16'h2142; weight[158] = 16'h9d3a; weight[159] = 16'hab33; weight[160] =
16'haf9b; weight[161] = 16'h2c0c; weight[162] = 16'h9cfb; weight[163] =
16'h26b0; weight[164] = 16'h2615; weight[165] = 16'h2d9a; weight[166] =
16'h2986; weight[167] = 16'hacd1; weight[168] = 16'hafba; weight[169] =
16'ha952; weight[170] = 16'h2e2e; weight[171] = 16'h25ff; weight[172] =
16'hac57; weight[173] = 16'h2693; weight[174] = 16'h2c2c; weight[175] =
16'hae57; weight[176] = 16'hb432; weight[177] = 16'h9a95; weight[178] =
16'ha044; weight[179] = 16'h9cc0; weight[180] = 16'had80; weight[181] =
16'hb166; weight[182] = 16'had51; weight[183] = 16'hb24e; weight[184] =
16'hb06d; weight[185] = 16'ha029; weight[186] = 16'h2d7c; weight[187] =
16'ha44a; weight[188] = 16'h0784; weight[189] = 16'ha8f0; weight[190] =
16'h28e1; weight[191] = 16'hadcf; weight[192] = 16'hae1e; weight[193] =
16'ha23d; weight[194] = 16'h26f8; weight[195] = 16'h2651; weight[196] =
16'h2080; weight[197] = 16'h29eb; weight[198] = 16'h247a; weight[199] =
16'hae97; weight[200] = 16'hadb6; weight[201] = 16'h22ef; weight[202] =
16'had7e; weight[203] = 16'h2677; weight[204] = 16'haab6; weight[205] =
16'ha297; weight[206] = 16'ha911; weight[207] = 16'hab18; weight[208] =
16'hacc5; weight[209] = 16'h2239; weight[210] = 16'ha279; weight[211] =
16'ha4ff; weight[212] = 16'h29e4; weight[213] = 16'h264b; weight[214] =
16'h91a9; weight[215] = 16'hac92; weight[216] = 16'ha4c4; weight[217] =
16'h2e10; weight[218] = 16'h2cf8; weight[219] = 16'h2823; weight[220] =
16'h2b09; weight[221] = 16'h2b32; weight[222] = 16'h9fbc; weight[223] =
16'h2953; weight[224] = 16'hac31; weight[225] = 16'h22f4; weight[226] =
16'h28b9; weight[227] = 16'h2db6; weight[228] = 16'h1c13; weight[229] =
16'h2590; weight[230] = 16'ha9a5; weight[231] = 16'h28b6; weight[232] =
16'ha966; weight[233] = 16'h3011; weight[234] = 16'h2b72; weight[235] =
16'h2f12; weight[236] = 16'h2cd7; weight[237] = 16'h2bbe; weight[238] =
16'h25cf; weight[239] = 16'h2b12; weight[240] = 16'habd5; weight[241] =
16'h299b; weight[242] = 16'h290c; weight[243] = 16'h31b4; weight[244] =
16'h25ef; weight[245] = 16'h2013; weight[246] = 16'h2908; weight[247] =
16'h293a; weight[248] = 16'hb072; weight[249] = 16'hb17e; weight[250] =
16'habc6; weight[251] = 16'h2c5c; weight[252] = 16'hb038; weight[253] =
16'hb185; weight[254] = 16'hb1fd; weight[255] = 16'hafc4; weight[256] =
16'hac9f; weight[257] = 16'h2dce; weight[258] = 16'h252e; weight[259] =
16'h329c; weight[260] = 16'h213f; weight[261] = 16'h21fd; weight[262] =
16'h223f; weight[263] = 16'ha41e; weight[264] = 16'haa1c; weight[265] =
16'h28fe; weight[266] = 16'h247c; weight[267] = 16'h297b; weight[268] =
16'h2878; weight[269] = 16'h2a86; weight[270] = 16'h20d2; weight[271] =
16'h2aa6; weight[272] = 16'had9d; weight[273] = 16'ha42a; weight[274] =
16'h1ddf; weight[275] = 16'h2fb7; weight[276] = 16'ha71a; weight[277] =
16'h25ba; weight[278] = 16'ha974; weight[279] = 16'ha46c; weight[280] =
16'haa92; weight[281] = 16'h2ca5; weight[282] = 16'h1cf1; weight[283] =
16'h29c6; weight[284] = 16'h27ea; weight[285] = 16'h2bb1; weight[286] =
16'h20b9; weight[287] = 16'h2828; weight[288] = 16'h9bbd; weight[289] =
16'h2135; weight[290] = 16'ha358; weight[291] = 16'ha9b5; weight[292] =
16'h2903; weight[293] = 16'h1cbd; weight[294] = 16'ha495; weight[295] =
16'h28e0; weight[296] = 16'h9c16; weight[297] = 16'had99; weight[298] =
16'haa51; weight[299] = 16'ha618; weight[300] = 16'ha57d; weight[301] =
16'haa74; weight[302] = 16'h2c99; weight[303] = 16'ha863; weight[304] =
16'h2866; weight[305] = 16'ha52d; weight[306] = 16'h9efa; weight[307] =
16'ha0ce; weight[308] = 16'h2893; weight[309] = 16'h2992; weight[310] =
16'h1f34; weight[311] = 16'h2553; weight[312] = 16'hac44; weight[313] =
16'h29ff; weight[314] = 16'h2078; weight[315] = 16'hb364; weight[316] =
16'h2948; weight[317] = 16'h25eb; weight[318] = 16'h16bc; weight[319] =
16'h24a2; weight[320] = 16'hab3c; weight[321] = 16'had56; weight[322] =
16'ha733; weight[323] = 16'haf34; weight[324] = 16'h2c08; weight[325] =
16'hae47; weight[326] = 16'h24ee; weight[327] = 16'hade6; weight[328] =
16'h279f; weight[329] = 16'haf72; weight[330] = 16'ha50e; weight[331] =
16'h2b14; weight[332] = 16'h1670; weight[333] = 16'h240f; weight[334] =
16'h9cf4; weight[335] = 16'ha688; weight[336] = 16'ha984; weight[337] =
16'h2899; weight[338] = 16'h283a; weight[339] = 16'haab3; weight[340] =
16'hab1e; weight[341] = 16'h25e5; weight[342] = 16'ha50e; weight[343] =
16'ha1ca; weight[344] = 16'h18d4; weight[345] = 16'h2985; weight[346] =
16'h297c; weight[347] = 16'h2800; weight[348] = 16'ha774; weight[349] =
16'h30ed; weight[350] = 16'ha76d; weight[351] = 16'h1545; weight[352] =
16'h29cc; weight[353] = 16'h2719; weight[354] = 16'h2db1; weight[355] =
16'h2921; weight[356] = 16'habdc; weight[357] = 16'h3091; weight[358] =
16'h9e15; weight[359] = 16'ha76d; weight[360] = 16'h257e; weight[361] =
16'h1d16; weight[362] = 16'h24f7; weight[363] = 16'h2516; weight[364] =
16'h2de9; weight[365] = 16'ha7a2; weight[366] = 16'h26c9; weight[367] =
16'h25d4; weight[368] = 16'h25fe; weight[369] = 16'hada5; weight[370] =
16'h1c82; weight[371] = 16'ha805; weight[372] = 16'h2564; weight[373] =
16'h27b1; weight[374] = 16'ha44e; weight[375] = 16'hb48f; weight[376] =
16'h2c5c; weight[377] = 16'had75; weight[378] = 16'h29a4; weight[379] =
16'ha7e9; weight[380] = 16'h3042; weight[381] = 16'h2377; weight[382] =
16'hac5b; weight[383] = 16'h3138; weight[384] = 16'ha61c; weight[385] =
16'hb03d; weight[386] = 16'ha668; weight[387] = 16'h92af; weight[388] =
16'h25f9; weight[389] = 16'h236b; weight[390] = 16'h2ddd; weight[391] =
16'hadd6; weight[392] = 16'ha552; weight[393] = 16'hacc1; weight[394] =
16'hb38f; weight[395] = 16'h2c80; weight[396] = 16'ha835; weight[397] =
16'h28f3; weight[398] = 16'ha6d5; weight[399] = 16'hb607; weight[400] =
16'h26aa; weight[401] = 16'hb1a2; weight[402] = 16'h2bc3; weight[403] =
16'ha8de; weight[404] = 16'h27c2; weight[405] = 16'h2cb2; weight[406] =
16'hb157; weight[407] = 16'h30ae; weight[408] = 16'h1178; weight[409] =
16'hb008; weight[410] = 16'h2ee0; weight[411] = 16'ha3d8; weight[412] =
16'ha88f; weight[413] = 16'hadd1; weight[414] = 16'h287a; weight[415] =
16'h3198; weight[416] = 16'h1cfa; weight[417] = 16'hb351; weight[418] =
16'ha2c1; weight[419] = 16'ha4c4; weight[420] = 16'hac69; weight[421] =
16'hb10c; weight[422] = 16'ha5b5; weight[423] = 16'h325f; weight[424] =
16'ha56e; weight[425] = 16'hb099; weight[426] = 16'h3002; weight[427] =
16'h228b; weight[428] = 16'ha1cc; weight[429] = 16'had2a; weight[430] =
16'h2061; weight[431] = 16'h35b4; weight[432] = 16'haaff; weight[433] =
16'h300b; weight[434] = 16'hab1d; weight[435] = 16'h2d66; weight[436] =
16'h329d; weight[437] = 16'h238d; weight[438] = 16'h9833; weight[439] =
16'haafc; weight[440] = 16'h1fa7; weight[441] = 16'h2971; weight[442] =
16'h20df; weight[443] = 16'h2c42; weight[444] = 16'h2d90; weight[445] =
16'h2e5a; weight[446] = 16'h289f; weight[447] = 16'h2825; weight[448] =
16'had18; weight[449] = 16'h2a4b; weight[450] = 16'h2588; weight[451] =
16'h2e73; weight[452] = 16'h9d0e; weight[453] = 16'h277a; weight[454] =
16'h1653; weight[455] = 16'ha1ab; weight[456] = 16'h200e; weight[457] =
16'h2e51; weight[458] = 16'ha924; weight[459] = 16'h2953; weight[460] =
16'h33a9; weight[461] = 16'h28a3; weight[462] = 16'h2382; weight[463] =
16'ha6f3; weight[464] = 16'h29a1; weight[465] = 16'ha898; weight[466] =
16'h2c18; weight[467] = 16'h1fde; weight[468] = 16'hb20b; weight[469] =
16'ha526; weight[470] = 16'ha9d2; weight[471] = 16'h2435; weight[472] =
16'h2705; weight[473] = 16'ha558; weight[474] = 16'h309d; weight[475] =
16'h2c18; weight[476] = 16'hb2a6; weight[477] = 16'h1a43; weight[478] =
16'ha754; weight[479] = 16'h2c53; weight[480] = 16'ha736; weight[481] =
16'h2b03; weight[482] = 16'ha674; weight[483] = 16'h211a; weight[484] =
16'h2939; weight[485] = 16'hab9c; weight[486] = 16'h2a93; weight[487] =
16'ha27b; weight[488] = 16'ha413; weight[489] = 16'h24e4; weight[490] =
16'h2c91; weight[491] = 16'h9a53; weight[492] = 16'haf36; weight[493] =
16'haa7e; weight[494] = 16'h2614; weight[495] = 16'h21ea; weight[496] =
16'ha3c3; weight[497] = 16'ha7d2; weight[498] = 16'h2c93; weight[499] =
16'h2856; weight[500] = 16'ha58e; weight[501] = 16'h189f; weight[502] =
16'ha4f1; weight[503] = 16'ha26e; weight[504] = 16'hb174; weight[505] =
16'ha9df; weight[506] = 16'hac27; weight[507] = 16'haa2d; weight[508] =
16'h284c; weight[509] = 16'ha5a8; weight[510] = 16'hac9e; weight[511] =
16'had61; weight[512] = 16'h2433; weight[513] = 16'h2bdc; weight[514] =
16'ha6de; weight[515] = 16'h28a5; weight[516] = 16'h2a42; weight[517] =
16'ha159; weight[518] = 16'h285e; weight[519] = 16'had2a; weight[520] =
16'ha220; weight[521] = 16'ha984; weight[522] = 16'ha37d; weight[523] =
16'ha83e; weight[524] = 16'ha87f; weight[525] = 16'h9c86; weight[526] =
16'h236b; weight[527] = 16'h8ca1; weight[528] = 16'hb13f; weight[529] =
16'hac1d; weight[530] = 16'ha615; weight[531] = 16'h2cad; weight[532] =
16'h2a9d; weight[533] = 16'h2a88; weight[534] = 16'ha208; weight[535] =
16'ha75c; weight[536] = 16'h1827; weight[537] = 16'h2c74; weight[538] =
16'ha8b0; weight[539] = 16'ha94a; weight[540] = 16'ha95c; weight[541] =
16'had39; weight[542] = 16'h2b86; weight[543] = 16'hae38; weight[544] =
16'h309d; weight[545] = 16'ha606; weight[546] = 16'h2a9c; weight[547] =
16'h2ccf; weight[548] = 16'hac28; weight[549] = 16'hac53; weight[550] =
16'h2d39; weight[551] = 16'h2805; weight[552] = 16'ha59d; weight[553] =
16'hac43; weight[554] = 16'h2603; weight[555] = 16'h28c2; weight[556] =
16'h27e1; weight[557] = 16'h2e48; weight[558] = 16'h1f11; weight[559] =
16'ha17e; weight[560] = 16'h2267; weight[561] = 16'h29ba; weight[562] =
16'ha969; weight[563] = 16'habaa; weight[564] = 16'ha0d8; weight[565] =
16'h2bba; weight[566] = 16'h2bbb; weight[567] = 16'h1f7f; weight[568] =
16'h2daf; weight[569] = 16'hac8c; weight[570] = 16'h26e1; weight[571] =
16'h1f08; weight[572] = 16'ha6eb; weight[573] = 16'h2362; weight[574] =
16'h2659; weight[575] = 16'h2802; weight[576] = 16'h30ac; weight[577] =
16'habd1; weight[578] = 16'ha637; weight[579] = 16'ha99b; weight[580] =
16'h2a89; weight[581] = 16'h193a; weight[582] = 16'ha51c; weight[583] =
16'h2fde; weight[584] = 16'h2e59; weight[585] = 16'hae16; weight[586] =
16'h26d6; weight[587] = 16'haf5e; weight[588] = 16'hacea; weight[589] =
16'ha9c5; weight[590] = 16'ha70c; weight[591] = 16'h29a2; weight[592] =
16'h29b4; weight[593] = 16'h25d6; weight[594] = 16'h26df; weight[595] =
16'hac37; weight[596] = 16'ha5c4; weight[597] = 16'h2def; weight[598] =
16'h26b2; weight[599] = 16'h2d4f; weight[600] = 16'h2a2b; weight[601] =
16'hac19; weight[602] = 16'haef5; weight[603] = 16'ha422; weight[604] =
16'h2f0d; weight[605] = 16'h2683; weight[606] = 16'h257c; weight[607] =
16'h2ef4; weight[608] = 16'h2c13; weight[609] = 16'haa70; weight[610] =
16'hae4d; weight[611] = 16'haa46; weight[612] = 16'hab07; weight[613] =
16'haf00; weight[614] = 16'ha9ed; weight[615] = 16'ha613; weight[616] =
16'h2bd8; weight[617] = 16'h292c; weight[618] = 16'hadab; weight[619] =
16'habcf; weight[620] = 16'h23a3; weight[621] = 16'h2d3f; weight[622] =
16'h2841; weight[623] = 16'h2af0; weight[624] = 16'h2829; weight[625] =
16'ha964; weight[626] = 16'h258a; weight[627] = 16'hae39; weight[628] =
16'ha7d0; weight[629] = 16'h2a99; weight[630] = 16'h278c; weight[631] =
16'h2eb9; weight[632] = 16'h2d62; weight[633] = 16'haf62; weight[634] =
16'h2826; weight[635] = 16'haecc; weight[636] = 16'ha08e; weight[637] =
16'ha758; weight[638] = 16'h9e07; weight[639] = 16'h300f; weight[640] =
16'h31b0; weight[641] = 16'ha240; weight[642] = 16'h9f1b; weight[643] =
16'ha47d; weight[644] = 16'h29cb; weight[645] = 16'h2c75; weight[646] =
16'h239f; weight[647] = 16'h2dc7; weight[648] = 16'ha1f4; weight[649] =
16'h26f1; weight[650] = 16'h2508; weight[651] = 16'hb338; weight[652] =
16'h2713; weight[653] = 16'h99f7; weight[654] = 16'h2922; weight[655] =
16'h28ea; weight[656] = 16'h2e7d; weight[657] = 16'ha9d1; weight[658] =
16'h2694; weight[659] = 16'hb0a9; weight[660] = 16'ha08d; weight[661] =
16'ha55f; weight[662] = 16'h287f; weight[663] = 16'ha395; weight[664] =
16'haa99; weight[665] = 16'h2365; weight[666] = 16'h251f; weight[667] =
16'hb1db; weight[668] = 16'h1968; weight[669] = 16'h2bdb; weight[670] =
16'h002c; weight[671] = 16'h28e2; weight[672] = 16'hab35; weight[673] =
16'hac2b; weight[674] = 16'h279e; weight[675] = 16'hae6d; weight[676] =
16'h939b; weight[677] = 16'h21bc; weight[678] = 16'ha919; weight[679] =
16'hab85; weight[680] = 16'h174d; weight[681] = 16'hadf7; weight[682] =
16'h1d97; weight[683] = 16'ha239; weight[684] = 16'had16; weight[685] =
16'haf10; weight[686] = 16'h288b; weight[687] = 16'h9675; weight[688] =
16'had8f; weight[689] = 16'haaf6; weight[690] = 16'h23b9; weight[691] =
16'haf7e; weight[692] = 16'h1094; weight[693] = 16'h1fe9; weight[694] =
16'ha706; weight[695] = 16'h28f7; weight[696] = 16'hab55; weight[697] =
16'h2ae7; weight[698] = 16'hacd5; weight[699] = 16'hb3ef; weight[700] =
16'h2c61; weight[701] = 16'h2867; weight[702] = 16'ha0ce; weight[703] =
16'ha83a; weight[704] = 16'h2eb1; weight[705] = 16'h279f; weight[706] =
16'ha3a5; weight[707] = 16'hb231; weight[708] = 16'h9c86; weight[709] =
16'ha2b0; weight[710] = 16'h208a; weight[711] = 16'ha5f5; weight[712] =
16'haa23; weight[713] = 16'h2c9f; weight[714] = 16'h2c9c; weight[715] =
16'hb3f2; weight[716] = 16'h2afe; weight[717] = 16'h1876; weight[718] =
16'h21c8; weight[719] = 16'h2da3; weight[720] = 16'h2b5c; weight[721] =
16'h2d49; weight[722] = 16'h2d7c; weight[723] = 16'ha500; weight[724] =
16'ha9db; weight[725] = 16'ha970; weight[726] = 16'h265f; weight[727] =
16'ha54f; weight[728] = 16'h2551; weight[729] = 16'h2954; weight[730] =
16'h3012; weight[731] = 16'ha9c7; weight[732] = 16'ha8dd; weight[733] =
16'hacbd; weight[734] = 16'h20cf; weight[735] = 16'h1e5a; weight[736] =
16'ha75c; weight[737] = 16'h1769; weight[738] = 16'h2fce; weight[739] =
16'h2a7d; weight[740] = 16'h140c; weight[741] = 16'ha626; weight[742] =
16'h27ed; weight[743] = 16'h2a40; weight[744] = 16'ha689; weight[745] =
16'h1f91; weight[746] = 16'h1fa5; weight[747] = 16'ha0b5; weight[748] =
16'h9e83; weight[749] = 16'ha4fa; weight[750] = 16'h26cd; weight[751] =
16'h1ed8; weight[752] = 16'ha839; weight[753] = 16'ha38e; weight[754] =
16'h27ae; weight[755] = 16'ha5bd; weight[756] = 16'habcf; weight[757] =
16'ha0da; weight[758] = 16'h1e42; weight[759] = 16'ha905; weight[760] =
16'ha515; weight[761] = 16'ha830; weight[762] = 16'h2772; weight[763] =
16'h1dba; weight[764] = 16'ha416; weight[765] = 16'h1d0d; weight[766] =
16'ha40c; weight[767] = 16'ha58e; weight[768] = 16'ha9e8; weight[769] =
16'h9488; weight[770] = 16'ha601; weight[771] = 16'had44; weight[772] =
16'hac56; weight[773] = 16'h275d; weight[774] = 16'h2add; weight[775] =
16'ha7b4; weight[776] = 16'hae71; weight[777] = 16'hae16; weight[778] =
16'ha89e; weight[779] = 16'hadbc; weight[780] = 16'hb09d; weight[781] =
16'h24ee; weight[782] = 16'h25ed; weight[783] = 16'hb03a; weight[784] =
16'ha605; weight[785] = 16'hada6; weight[786] = 16'haeb2; weight[787] =
16'h9df5; weight[788] = 16'ha494; weight[789] = 16'h2b13; weight[790] =
16'h2a1f; weight[791] = 16'ha016; weight[792] = 16'h2d23; weight[793] =
16'h32a6; weight[794] = 16'h2ed6; weight[795] = 16'h214b; weight[796] =
16'h20a2; weight[797] = 16'h92be; weight[798] = 16'h283d; weight[799] =
16'h25e4; weight[800] = 16'h2a85; weight[801] = 16'h34dd; weight[802] =
16'h3007; weight[803] = 16'ha7b6; weight[804] = 16'h22ad; weight[805] =
16'h2109; weight[806] = 16'ha7cd; weight[807] = 16'hac30; weight[808] =
16'h2982; weight[809] = 16'h3346; weight[810] = 16'h2fcf; weight[811] =
16'h17c2; weight[812] = 16'h26d5; weight[813] = 16'h1c03; weight[814] =
16'habd6; weight[815] = 16'ha5c8; weight[816] = 16'h26a6; weight[817] =
16'h1c9c; weight[818] = 16'h287a; weight[819] = 16'ha453; weight[820] =
16'ha742; weight[821] = 16'ha64c; weight[822] = 16'h21c3; weight[823] =
16'h2c0f; weight[824] = 16'ha951; weight[825] = 16'h2c3e; weight[826] =
16'hafa8; weight[827] = 16'h9ca6; weight[828] = 16'haa12; weight[829] =
16'h20e2; weight[830] = 16'ha922; weight[831] = 16'h2d8d; weight[832] =
16'h2526; weight[833] = 16'h1e2a; weight[834] = 16'haa66; weight[835] =
16'ha620; weight[836] = 16'ha94d; weight[837] = 16'h2988; weight[838] =
16'h271d; weight[839] = 16'h2b5d; weight[840] = 16'h29a5; weight[841] =
16'hae38; weight[842] = 16'had12; weight[843] = 16'h2bb5; weight[844] =
16'ha778; weight[845] = 16'h259a; weight[846] = 16'h2757; weight[847] =
16'h9f2f; weight[848] = 16'ha473; weight[849] = 16'hb4d1; weight[850] =
16'hb084; weight[851] = 16'ha652; weight[852] = 16'had15; weight[853] =
16'h22fb; weight[854] = 16'haad8; weight[855] = 16'haf0c; weight[856] =
16'h28fb; weight[857] = 16'hb0a6; weight[858] = 16'hb109; weight[859] =
16'h2618; weight[860] = 16'ha402; weight[861] = 16'h2d0e; weight[862] =
16'h2aa0; weight[863] = 16'h9e53; weight[864] = 16'h2c82; weight[865] =
16'h9cc9; weight[866] = 16'h2ab4; weight[867] = 16'ha4d0; weight[868] =
16'h28bb; weight[869] = 16'h2fec; weight[870] = 16'h2603; weight[871] =
16'ha112; weight[872] = 16'hac6f; weight[873] = 16'haaea; weight[874] =
16'h1e69; weight[875] = 16'hb04e; weight[876] = 16'hb116; weight[877] =
16'haad0; weight[878] = 16'hacdb; weight[879] = 16'h0fd9; weight[880] =
16'hae4b; weight[881] = 16'ha5a6; weight[882] = 16'h272c; weight[883] =
16'h2d5c; weight[884] = 16'h27fb; weight[885] = 16'h2671; weight[886] =
16'h1789; weight[887] = 16'h2148; weight[888] = 16'ha856; weight[889] =
16'h1afd; weight[890] = 16'h260e; weight[891] = 16'ha3f4; weight[892] =
16'h1ffb; weight[893] = 16'ha2da; weight[894] = 16'ha07b; weight[895] =
16'ha670; weight[896] = 16'h2201; weight[897] = 16'h24ed; weight[898] =
16'haef8; weight[899] = 16'had4a; weight[900] = 16'h2eb6; weight[901] =
16'haf27; weight[902] = 16'ha0e8; weight[903] = 16'h2c1d; weight[904] =
16'h20ee; weight[905] = 16'h9490; weight[906] = 16'had88; weight[907] =
16'h2b29; weight[908] = 16'h2be9; weight[909] = 16'ha1a1; weight[910] =
16'hab45; weight[911] = 16'haf06; weight[912] = 16'had87; weight[913] =
16'ha33f; weight[914] = 16'h2ad1; weight[915] = 16'h2712; weight[916] =
16'ha615; weight[917] = 16'h2ffc; weight[918] = 16'h2eeb; weight[919] =
16'h2e5a; weight[920] = 16'ha585; weight[921] = 16'ha1b0; weight[922] =
16'ha570; weight[923] = 16'hb149; weight[924] = 16'hb13d; weight[925] =
16'habce; weight[926] = 16'h2ca7; weight[927] = 16'ha670; weight[928] =
16'h2a16; weight[929] = 16'h1ded; weight[930] = 16'ha891; weight[931] =
16'ha8de; weight[932] = 16'haa7f; weight[933] = 16'h2f13; weight[934] =
16'h2b31; weight[935] = 16'ha422; weight[936] = 16'h9fe7; weight[937] =
16'ha803; weight[938] = 16'ha3d7; weight[939] = 16'h2cba; weight[940] =
16'h27e8; weight[941] = 16'h9f6a; weight[942] = 16'ha088; weight[943] =
16'h30d9; weight[944] = 16'h280d; weight[945] = 16'h248d; weight[946] =
16'h27db; weight[947] = 16'hae09; weight[948] = 16'h31cb; weight[949] =
16'haab6; weight[950] = 16'h2890; weight[951] = 16'hb4d0; weight[952] =
16'ha457; weight[953] = 16'h24b4; weight[954] = 16'h262e; weight[955] =
16'h29b1; weight[956] = 16'h16d1; weight[957] = 16'hac5b; weight[958] =
16'hb030; weight[959] = 16'hac07; weight[960] = 16'hb226; weight[961] =
16'hb12d; weight[962] = 16'ha7a9; weight[963] = 16'hafc7; weight[964] =
16'ha9ac; weight[965] = 16'haca2; weight[966] = 16'hb088; weight[967] =
16'h30db; weight[968] = 16'h2e68; weight[969] = 16'h34c1; weight[970] =
16'ha91f; weight[971] = 16'h343b; weight[972] = 16'h3295; weight[973] =
16'h32eb; weight[974] = 16'h330f; weight[975] = 16'ha540; weight[976] =
16'hb040; weight[977] = 16'h2425; weight[978] = 16'hb0fd; weight[979] =
16'ha794; weight[980] = 16'ha7df; weight[981] = 16'ha4a3; weight[982] =
16'hb393; weight[983] = 16'h2274; weight[984] = 16'h06fe; weight[985] =
16'h21a3; weight[986] = 16'h3011; weight[987] = 16'h296a; weight[988] =
16'haf55; weight[989] = 16'had8b; weight[990] = 16'hb011; weight[991] =
16'h2f49; weight[992] = 16'h2976; weight[993] = 16'hae03; weight[994] =
16'h2c02; weight[995] = 16'hac11; weight[996] = 16'haaae; weight[997] =
16'h2d41; weight[998] = 16'h2771; weight[999] = 16'ha8b1; weight[1000] = 16'h2a5e; weight[1001] = 16'h2a55; weight[1002] = 16'h2119; weight[1003] = 16'h2a80; weight[1004] = 16'hac11; weight[1005] = 16'h15ab; weight[1006] = 16'h23e5; weight[1007] = 16'h2e49; weight[1008] = 16'h26ea; weight[1009] = 16'h2e10; weight[1010] = 16'hac52; weight[1011] = 16'h2965; weight[1012] = 16'h9826; weight[1013] = 16'h298e; weight[1014] = 16'h9d94; weight[1015] = 16'h252d; weight[1016] = 16'h2dc3; weight[1017] = 16'h3085; weight[1018] = 16'hb2cf; weight[1019] = 16'h31b7; weight[1020] = 16'h22b0; weight[1021] = 16'ha92b; weight[1022] = 16'hac87; weight[1023] =
16'ha530; weight[1024] = 16'h2974; weight[1025] = 16'h2a84; weight[1026] = 16'habac; weight[1027] = 16'h2cba; weight[1028] = 16'ha3b2; weight[1029] = 16'h2707; weight[1030] = 16'h2753; weight[1031] = 16'h2193; weight[1032] = 16'ha9b2; weight[1033] = 16'h9c59; weight[1034] = 16'had93; weight[1035] = 16'h2bff; weight[1036] = 16'h1d86; weight[1037] = 16'h9915;
weight[1038] = 16'h25a7; weight[1039] = 16'h2bd8; weight[1040] = 16'h2aee; weight[1041] = 16'hae1a; weight[1042] = 16'hb04d; weight[1043] = 16'ha6dd; weight[1044] = 16'h2c71; weight[1045] = 16'ha137; weight[1046] = 16'h26a2; weight[1047] = 16'h25f4; weight[1048] = 16'h1348; weight[1049]
= 16'h2758; weight[1050] = 16'haf1c; weight[1051] = 16'h13d5; weight[1052] = 16'h2ca3; weight[1053] = 16'h2612; weight[1054] = 16'h9caa; weight[1055] = 16'habf9; weight[1056] = 16'ha8dd; weight[1057] = 16'ha687; weight[1058] = 16'h2e1a; weight[1059] = 16'ha6d0; weight[1060] = 16'ha5d9; weight[1061] = 16'ha4b6; weight[1062] = 16'h2493; weight[1063] = 16'h2866; weight[1064] = 16'ha9dd; weight[1065] = 16'haddf; weight[1066] = 16'h3316; weight[1067] = 16'hb1ce; weight[1068] = 16'hae2f; weight[1069] = 16'h999c; weight[1070] = 16'h2b48; weight[1071] = 16'h2854; weight[1072] = 16'h2add; weight[1073] = 16'ha1e2; weight[1074] = 16'h2a96; weight[1075] = 16'ha9b6; weight[1076] = 16'ha474; weight[1077] = 16'haa64; weight[1078] = 16'haa2a; weight[1079] = 16'hac22; weight[1080] = 16'hadd2; weight[1081] = 16'h9459; weight[1082] = 16'ha527; weight[1083] = 16'ha7b4; weight[1084] = 16'h2529; weight[1085] = 16'h2c58; weight[1086] = 16'h299c; weight[1087] = 16'ha1e8; weight[1088] = 16'hb8b4; weight[1089] = 16'ha785; weight[1090] = 16'h20e2; weight[1091] = 16'had11; weight[1092] = 16'h18bb; weight[1093] = 16'ha555; weight[1094] = 16'hb33e; weight[1095] =
16'h2774; weight[1096] = 16'h28c1; weight[1097] = 16'h0e17; weight[1098] = 16'ha07f; weight[1099] = 16'ha040; weight[1100] = 16'h2920; weight[1101] = 16'h290d; weight[1102] = 16'h242d; weight[1103] = 16'h25be; weight[1104] = 16'ha097; weight[1105] = 16'ha64e; weight[1106] = 16'hac79; weight[1107] = 16'h21f1; weight[1108] = 16'ha202; weight[1109] = 16'h1594;
weight[1110] = 16'h1b6b; weight[1111] = 16'h1e7b; weight[1112] = 16'ha695; weight[1113] = 16'h1737; weight[1114] = 16'h1c3a; weight[1115] = 16'h2dd9; weight[1116] = 16'ha11d; weight[1117] = 16'h2a2b; weight[1118] = 16'ha7de; weight[1119] = 16'h2677; weight[1120] = 16'hac8c; weight[1121]
= 16'ha811; weight[1122] = 16'h1eb7; weight[1123] = 16'had35; weight[1124] = 16'h1e13; weight[1125] = 16'h9872; weight[1126] = 16'h28da; weight[1127] = 16'h9caa; weight[1128] = 16'h2e19; weight[1129] = 16'h9de5; weight[1130] = 16'ha946; weight[1131] = 16'h9ae5; weight[1132] = 16'ha5f9; weight[1133] = 16'hada0; weight[1134] = 16'ha7f8; weight[1135] = 16'h281a; weight[1136] = 16'h36bc; weight[1137] = 16'h2d25; weight[1138] = 16'ha85f; weight[1139] = 16'h2c82; weight[1140] = 16'ha5ba; weight[1141] = 16'h2499; weight[1142] = 16'h30a2; weight[1143] = 16'haa7d; weight[1144] = 16'h2c11; weight[1145] = 16'h241f; weight[1146] = 16'h23f4; weight[1147] = 16'ha6dd; weight[1148] = 16'ha9b4; weight[1149] = 16'ha374; weight[1150] = 16'h24a8; weight[1151] = 16'ha500;

	end
`endif
`ifdef SACC
	reg [169*16-1:0] avepooldata;
	initial begin
		avepooldata = {16'h3757, 16'h39da, 16'h3b67, 16'h3376, 16'h3bb5, 16'h30da, 16'h3b8a, 16'h2675, 16'h3454, 16'h2d3e, 16'h39d1, 16'h3614, 16'h36dd,
	16'h304e, 16'h3023, 16'h3b02, 16'h3367, 16'h3b9d, 16'h32ff, 16'h387e, 16'h384d, 16'h3812, 16'h3bad, 16'h3587, 16'h33f5, 16'h3ab1,
	16'h3945, 16'h3625, 16'h2f8f, 16'h39de, 16'h367c, 16'h287c, 16'h354f, 16'h2d21, 16'h39a8, 16'h382e, 16'h3b5c, 16'h3ba0, 16'h39cd,
	16'h3a0c, 16'h2e91, 16'h38cb, 16'h2bc9, 16'h3872, 16'h3173, 16'h37b0, 16'h32da, 16'h3b5a, 16'h380e, 16'h3892, 16'h3988, 16'h390d,
	16'h38e9, 16'h3a7c, 16'h3a78, 16'h3a50, 16'h3894, 16'h397d, 16'h314d, 16'h2c73, 16'h304c, 16'h3774, 16'h36ca, 16'h3512, 16'h3b17,
	16'h363f, 16'h3721, 16'h3489, 16'h2fe5, 16'h34c6, 16'h3aaf, 16'h37b1, 16'h38e3, 16'h36e3, 16'h3942, 16'h3bbe, 16'h39ac, 16'h3873,
	16'h37c1, 16'h340b, 16'h3b26, 16'h3b70, 16'h372c, 16'h36f3, 16'h3bd5, 16'h3a3a, 16'h339e, 16'h3821, 16'h33f5, 16'h3858, 16'h3bf0,
	16'h3beb, 16'h3b73, 16'h3a1c, 16'h3a83, 16'h3bb2, 16'h3808, 16'h39c7, 16'h3b72, 16'h39cf, 16'h2a93, 16'h3402, 16'h39d8, 16'h3974,
	16'h3483, 16'h3b46, 16'h3af9, 16'h38ad, 16'h3933, 16'h30de, 16'h305e, 16'h2fdb, 16'h3ad9, 16'h3ad2, 16'h39fa, 16'h2ae8, 16'h32b6,
	16'h3596, 16'h3b5e, 16'h329c, 16'h2da6, 16'h3a5a, 16'h3562, 16'h3a02, 16'h3a38, 16'h354e, 16'h3b19, 16'h3976, 16'h383c, 16'h29d8,
	16'h3a29, 16'h3a08, 16'h3301, 16'h386f, 16'h2a75, 16'h37cf, 16'h3267, 16'h30e1, 16'h3967, 16'h388a, 16'h397b, 16'h3ab4, 16'h3999,
	16'h3899, 16'h378f, 16'h394b, 16'h3554, 16'h3723, 16'h3880, 16'h327a, 16'h3a9b, 16'h383c, 16'h3936, 16'h387d, 16'h34c5, 16'h3782,
	16'h3a3f, 16'h3b8c, 16'h3156, 16'h3ba7, 16'h3b97, 16'h2e65, 16'h3194, 16'h32d6, 16'h3572, 16'h3889, 16'h3aa1, 16'h36d4, 16'h2cc5}; //16'h558f, 16'h3836
	end
`endif
`ifdef SCMP
	reg [127:0] maxpooldata[0:18];
	initial begin
		maxpooldata[0] = 128'h47505861000000000000000000004167;
		maxpooldata[1] = 128'h49045930000000000000000000004D86;
		maxpooldata[2] = 128'h48A659B938184A1E0000477B45E24C9A;
		maxpooldata[3] = 128'h4D10591D0000450D00000000482C0000;
		maxpooldata[4] = 128'h4B67592E00004B7C0000000048E20000;
		maxpooldata[5] = 128'h0000593B4269000000004A184B154B47;
		maxpooldata[6] = 128'h4D2F595D000043F1000000004CBD0000;
		maxpooldata[7] = 128'h00005900000000000000000000000000;
		maxpooldata[8] = 128'h3F7858D341E500000000484043624C92;
	end
`endif

engine engine_(
	.clk					(clk),
//Control signals csb->engine
	.rst					(rst),
	.engine_valid			(engine_valid),
	.op_type				(op_type),
	.stride					(stride),
	.stride2				(stride2),
	.kernel					(kernel),
	.kernel_size			(kernel_size),
	.i_channel				(i_channel),
	.o_channel				(o_channel),
	.i_side					(i_side),
	.o_side					(o_side),
	.bias					(bias),
//Response signals engine->csb
	.gemm_finish			(gemm_finish),
//Command path engine->dma
	.output_en		(output_en),
	.d_ram_read_addr		(d_ram_read_addr),
	.w_ram_read_addr		(w_ram_read_addr),
//Data path dma->engine
	.input_data			(input_data),
	.input_weig			(input_weig),
	.output_data			(output_data)
);

always #5 clk = ~clk;
always @(posedge clk) begin
	if(gemm_finish) engine_valid <= 0; // pull down engine_valid after the whole op is done
end

initial begin
    rst = 1;
    clk = 0;
    engine_valid = 0;
    op_type = 0; stride = 0; stride2 = 0;
	kernel = 0; kernel_size = 0; i_channel = 0; o_channel = 0; i_side = 0; o_side = 0; 
	input_data = 'd0;
	input_weig = 'd0;
	bias = 16'h0000;
    #20 rst = 1;
    #10 rst = 0;
`ifdef CMAC
	//3x3
    #100 op_type = 1; stride = 1; stride2 = 3;
		kernel = 3; kernel_size = 9; i_channel = 16; o_channel = 64; i_side = 56; o_side = 56; bias = 16'hAC88;//16'hA35C;
	//1x1
	// #100 op_type = 1; stride = 1; stride2 = 1;
		// kernel = 1; kernel_size = 1; i_channel = 64; o_channel = 16; i_side = 56; o_side = 56; bias = 16'hAC88;
`endif
`ifdef SCMP
	#100 op_type = 2; stride = 2; stride2 = 6;
		kernel = 3; kernel_size = 9; i_channel = 64; o_channel = 64; i_side = 113; o_side = 56; bias = 16'h0000;
`endif
`ifdef SACC
	#100 op_type = 3; stride = 1; 
		kernel = 13; kernel_size = 169; i_channel = 1000; o_channel = 1000; i_side = 13; o_side = 1; bias = 16'h0000;
`endif
    #10 engine_valid = 1;
	//#3000 rst = 1;
	//#20 rst = 0;
	//#20 engine_valid = 1;
end

always @(posedge clk) begin
`ifdef CMAC
	input_data <= {data[d_ram_read_addr*8+7], data[d_ram_read_addr*8+6], data[d_ram_read_addr*8+5], data[d_ram_read_addr*8+4], data[d_ram_read_addr*8+3], data[d_ram_read_addr*8+2], data[d_ram_read_addr*8+1], data[d_ram_read_addr*8+0]};
	input_weig <= {weight[w_ram_read_addr*8+7], weight[w_ram_read_addr*8+6], weight[w_ram_read_addr*8+5], weight[w_ram_read_addr*8+4], weight[w_ram_read_addr*8+3], weight[w_ram_read_addr*8+2], weight[w_ram_read_addr*8+1], weight[w_ram_read_addr*8+0]};
`endif
`ifdef SCMP
	input_data <= maxpooldata[d_ram_read_addr];
`endif
`ifdef SACC
	input_data <= {16{avepooldata[d_ram_read_addr*16 +: 16]}};
`endif
end
endmodule