module dma(
    input clk,
    input rst_n,
    input addr,
    input dma_ready,
    output dma_valid,
    output [127:0] data
);


endmodule