`timescale 1ns/1ps
`define CMAC
// `define SACC
// `define SCMP

module engine_tb;

reg 		clk;
//Control signals csb->engine
reg 		rst;
reg 		engine_valid;
reg [2:0] 	op_type;
reg	[3:0]	stride;
reg [15:0]  stride2;
reg [7:0]  	kernel;
reg [7:0]	kernel_size;
reg [15:0]  i_channel;
reg [15:0]  o_channel;
reg [7:0]	i_side;
reg [7:0]   o_side;
reg	[15:0]  bias;
//Response signals engine->csb
wire		gemm_finish;
wire 		engine_ready;
//Command path engine->dma
wire        dma_p0_writes_en;
wire        dma_p2_reads_en;
wire        dma_p3_reads_en;
//Data path dma->engine
reg [15:0] 	dma_p2_ob_data;
reg [15:0] 	dma_p3_ob_data;
reg 		dma_p2_ob_we;
reg 		dma_p3_ob_we;
//Data path engine->dma
wire [15:0]	dma_p0_ib_data;

`ifdef CMAC
	reg [15:0] data [0:216];
	reg [15:0] weight [0:72];
	initial begin
	data[0] = 16'hce83; data[1] = 16'h4f98; data[2] = 16'h4e17; data[3] = 16'h0000; 
	data[4] = 16'h0000; data[5] = 16'h0000; data[6] = 16'h0000; data[7] = 16'h0000; 
	data[8] = 16'hce24; data[9] = 16'h5087; data[10] = 16'h4F8D; data[11] = 16'h0000; 
	data[12] = 16'h0000; data[13] = 16'h0000; data[14] = 16'h0000; data[15] = 16'h0000; 
	data[16] = 16'hCCEF; data[17] = 16'h51FB; data[18] = 16'h50DE; data[19] = 16'h0000;
	data[20] = 16'h0000; data[21] = 16'h0000; data[22] = 16'h0000; data[23] = 16'h0000;

	data[24] = 16'hCDE5; data[25] = 16'h5087; data[26] = 16'h4F10; data[27] = 16'h0000; 
	data[28] = 16'h0000; data[29] = 16'h0000; data[30] = 16'h0000; data[31] = 16'h0000; 
	data[32] = 16'hCFEB; data[33] = 16'h4FA7; data[34] = 16'h4DA9; data[35] = 16'h0000; 
	data[36] = 16'h0000; data[37] = 16'h0000; data[38] = 16'h0000; data[39] = 16'h0000;
	data[40] = 16'hD035; data[41] = 16'h5050; data[42] = 16'h4E61; data[43] = 16'h0000; 
	data[44] = 16'h0000; data[45] = 16'h0000; data[46] = 16'h0000; data[47] = 16'h0000;

	data[48] = 16'hD0A0; data[49] = 16'h4E32; data[50] = 16'h4C33; data[51] = 16'h0000; 
	data[52] = 16'h0000; data[53] = 16'h0000; data[54] = 16'h0000; data[55] = 16'h0000; 
	data[56] = 16'hD151; data[57] = 16'h4D6D; data[58] = 16'h49E7; data[59] = 16'h0000;
	data[60] = 16'h0000; data[61] = 16'h0000; data[62] = 16'h0000; data[63] = 16'h0000; 
	data[64] = 16'hD157; data[65] = 16'h4E9C; data[66] = 16'h4BC3; data[67] = 16'h0000; 
	data[68] = 16'h0000; data[69] = 16'h0000; data[70] = 16'h0000; data[71] = 16'h0000; 
	
	data[72] = 16'hd2b2; data[73] = 16'h4bef; data[74] = 16'h405e; data[75] = 16'h0000; 
	data[76] = 16'h0000; data[77] = 16'h0000; data[78] = 16'h0000; data[79] = 16'h0000; 
	data[80] = 16'hd1fc; data[81] = 16'h4d8b; data[82] = 16'h482d; data[83] = 16'h0000;
	data[84] = 16'h0000; data[85] = 16'h0000; data[86] = 16'h0000; data[87] = 16'h0000; 
	data[88] = 16'hd1db; data[89] = 16'h4e52; data[90] = 16'h49b4; data[91] = 16'h0000;
	data[92] = 16'h0000; data[93] = 16'h0000; data[94] = 16'h0000; data[95] = 16'h0000; 

	data[96] = 16'hd37e; data[97] = 16'h4bba; data[98] = 16'h387c; data[99] = 16'h0000;
	data[100] = 16'h0000; data[101] = 16'h0000; data[102] = 16'h0000; data[103] = 16'h0000; 
	data[104] = 16'hd34c; data[105] = 16'h4c67; data[106] = 16'h414e; data[107] = 16'h0000;
	data[108] = 16'h0000; data[109] = 16'h0000; data[110] = 16'h0000; data[111] = 16'h0000; 
	data[112] = 16'hd2d5; data[113] = 16'h4cad; data[114] = 16'h44ab; data[115] = 16'h0000;
	data[116] = 16'h0000; data[117] = 16'h0000; data[118] = 16'h0000; data[119] = 16'h0000; 

	data[120] = 16'hd43b; data[121] = 16'h480b; data[122] = 16'hc7ca; data[123] = 16'h0000;
	data[124] = 16'h0000; data[125] = 16'h0000; data[126] = 16'h0000; data[127] = 16'h0000; 
	data[128] = 16'hd453; data[129] = 16'h472b; data[130] = 16'hc863; data[131] = 16'h0000;
	data[132] = 16'h0000; data[133] = 16'h0000; data[134] = 16'h0000; data[135] = 16'h0000; 
	data[136] = 16'hd30c; data[137] = 16'h4c7e; data[138] = 16'h4030; data[139] = 16'h0000;
	data[140] = 16'h0000; data[141] = 16'h0000; data[142] = 16'h0000; data[143] = 16'h0000;

	data[144] = 16'hd29a; data[145] = 16'h4c60; data[146] = 16'h40ea; data[147] = 16'h0000;
	data[148] = 16'h0000; data[149] = 16'h0000; data[150] = 16'h0000; data[151] = 16'h0000;
	data[152] = 16'hd2ce; data[153] = 16'h4b51; data[154] = 16'hb765; data[155] = 16'h0000;
	data[156] = 16'h0000; data[157] = 16'h0000; data[158] = 16'h0000; data[159] = 16'h0000;
	data[160] = 16'hd0e5; data[161] = 16'h4efb; data[162] = 16'h4988; data[163] = 16'h0000;
	data[164] = 16'h0000; data[165] = 16'h0000; data[166] = 16'h0000; data[167] = 16'h0000;

	data[168] = 16'hd012; data[169] = 16'h5035; data[170] = 16'h4cad; data[171] = 16'h0000;
	data[172] = 16'h0000; data[173] = 16'h0000; data[174] = 16'h0000; data[175] = 16'h0000;
	data[176] = 16'hd05e; data[177] = 16'h4f76; data[178] = 16'h4bdc; data[179] = 16'h0000;
	data[180] = 16'h0000; data[181] = 16'h0000; data[182] = 16'h0000; data[183] = 16'h0000;
	data[184] = 16'hcfee; data[185] = 16'h4ffd; data[186] = 16'h4b86; data[187] = 16'h0000;
	data[188] = 16'h0000; data[189] = 16'h0000; data[190] = 16'h0000; data[191] = 16'h0000;

	data[192] = 16'hd041; data[193] = 16'h4ff3; data[194] = 16'h4c36; data[195] = 16'h0000;
	data[196] = 16'h0000; data[197] = 16'h0000; data[198] = 16'h0000; data[199] = 16'h0000;
	data[200] = 16'hd11b; data[201] = 16'h4de2; data[202] = 16'h48c0; data[203] = 16'h0000;
	data[204] = 16'h0000; data[205] = 16'h0000; data[206] = 16'h0000; data[207] = 16'h0000;
	data[208] = 16'hd1a2; data[209] = 16'h4c5c; data[210] = 16'h4237; data[211] = 16'h0000;
	data[212] = 16'h0000; data[213] = 16'h0000; data[214] = 16'h0000; data[215] = 16'h0000;

	weight[0] = 16'h341E; weight[1] = 16'h3867; weight[2] = 16'h3509; weight[3] = 16'h0000;
	weight[4] = 16'h0000; weight[5] = 16'h0000; weight[6] = 16'h0000; weight[7] = 16'h0000;
	weight[8] = 16'hAE6E; weight[9] = 16'hB0BF;	weight[10] = 16'hB0F7; weight[11] = 16'h0000;
	weight[12] = 16'h0000; weight[13] = 16'h0000; weight[14] = 16'h0000; weight[15] = 16'h0000;
	weight[16] = 16'hAC84; weight[17] = 16'hB2B4; weight[18] = 16'hAF54; weight[19] = 16'h0000;
	weight[20] = 16'h0000; weight[21] = 16'h0000; weight[22] = 16'h0000; weight[23] = 16'h0000;

	weight[24] = 16'h35C0; weight[25] = 16'h396D; weight[26] = 16'h36E1; weight[27] = 16'h0000;
	weight[28] = 16'h0000; weight[29] = 16'h0000; weight[30] = 16'h0000; weight[31] = 16'h0000;
	weight[32] = 16'hB10F; weight[33] = 16'hB456; weight[34] = 16'hB2C4; weight[35] = 16'h0000;
	weight[36] = 16'h0000; weight[37] = 16'h0000; weight[38] = 16'h0000; weight[39] = 16'h0000;
	weight[40] = 16'hB209; weight[41] = 16'hB76D; weight[42] = 16'hB3F0; weight[43] = 16'h0000;
	weight[44] = 16'h0000; weight[45] = 16'h0000; weight[46] = 16'h0000; weight[47] = 16'h0000;

	weight[48] = 16'h3282; weight[49] = 16'h376F; weight[50] = 16'h3504; weight[51] = 16'h0000;
	weight[52] = 16'h0000; weight[53] = 16'h0000; weight[54] = 16'h0000; weight[55] = 16'h0000;
	weight[56] = 16'hAE46; weight[57] = 16'hB1E7; weight[58] = 16'hACF0; weight[59] = 16'h0000;
	weight[60] = 16'h0000; weight[61] = 16'h0000; weight[62] = 16'h0000; weight[63] = 16'h0000;
	weight[64] = 16'hB249; weight[65] = 16'hB72B; weight[66] = 16'hB338; weight[67] = 16'h0000;
	weight[68] = 16'h0000; weight[69] = 16'h0000; weight[70] = 16'h0000; weight[71] = 16'h0000;
/*

d1f000004d030000451a00000000000000000000000000000000000000000000
d2fa000049270000c49500000000000000000000000000000000000000000000
d3d100003e840000ca3400000000000000000000000000000000000000000000
d374000048f00000c43800000000000000000000000000000000000000000000
d3920000489d0000c4ed00000000000000000000000000000000000000000000
d311000048690000c45d00000000000000000000000000000000000000000000
d440000044490000c8d600000000000000000000000000000000000000000000
d33a00004b8800003c3900000000000000000000000000000000000000000000
d2c900004bb500003e3400000000000000000000000000000000000000000000
d47c000046d90000c7f000000000000000000000000000000000000000000000
d3e100004b430000b52700000000000000000000000000000000000000000000
d40d000049500000c43800000000000000000000000000000000000000000000
d469000045df0000c88a00000000000000000000000000000000000000000000
d30300004d280000459d00000000000000000000000000000000000000000000
d28b00004d680000476a00000000000000000000000000000000000000000000
d32c0000492b0000c49d00000000000000000000000000000000000000000000
d0e000004f4f00004b1e00000000000000000000000000000000000000000000
cf48000050a000004dbe00000000000000000000000000000000000000000000
d1ce00004c0e0000401d00000000000000000000000000000000000000000000
cedc0000504500004cfd00000000000000000000000000000000000000000000
cd420000510400004e8800000000000000000000000000000000000000000000
d18d00004cc0000045d000000000000000000000000000000000000000000000
ce8a0000506100004da400000000000000000000000000000000000000000000
cc7c0000510500004ebe00000000000000000000000000000000000000000000
d1a500004d3d000047fd00000000000000000000000000000000000000000000
cef90000507a00004dc200000000000000000000000000000000000000000000
cec100004fa200004c6200000000000000000000000000000000000000000000
d1ad00004d5a0000483900000000000000000000000000000000000000000000
d14d00004dae000048db00000000000000000000000000000000000000000000
d25c000049300000c2ba00000000000000000000000000000000000000000000
d20b00004d8a0000483900000000000000000000000000000000000000000000
d1e100004cf8000046db00000000000000000000000000000000000000000000
d3a7000041610000c9a500000000000000000000000000000000000000000000
d14400004f6a00004bd900000000000000000000000000000000000000000000
d1dd00004dab0000487800000000000000000000000000000000000000000000
d35f000046f70000c7bd00000000000000000000000000000000000000000000
d09300004fe800004c9800000000000000000000000000000000000000000000
d1ac00004db4000048c200000000000000000000000000000000000000000000
d1e700004c730000431500000000000000000000000000000000000000000000
d13800004c85000045d200000000000000000000000000000000000000000000
d3c50000bf5c0000cb1300000000000000000000000000000000000000000000
d35300003ac90000c9e000000000000000000000000000000000000000000000
d10900004a3c00003cbf00000000000000000000000000000000000000000000
d2a600003d730000c8fb00000000000000000000000000000000000000000000
d11400004afa0000414400000000000000000000000000000000000000000000
d07800004c200000458700000000000000000000000000000000000000000000
d01100004d32000048e300000000000000000000000000000000000000000000
ccd40000504100004dc100000000000000000000000000000000000000000000
cdfc00004e6b00004bae00000000000000000000000000000000000000000000
cdad00004ed400004c3e00000000000000000000000000000000000000000000
ccdb00004fa600004d1000000000000000000000000000000000000000000000
ce1900004ceb0000492b00000000000000000000000000000000000000000000
ce1000004d0c0000496a00000000000000000000000000000000000000000000
cdd600004d47000049df00000000000000000000000000000000000000000000
cd9d00004c90000048a200000000000000000000000000000000000000000000
cc9c00004da800004acf00000000000000000000000000000000000000000000
cbe900004e9f00004c5e00000000000000000000000000000000000000000000
cb9e00004f1e00004cb700000000000000000000000000000000000000000000
c8df0000504b00004e2d00000000000000000000000000000000000000000000
c4ef000050d500004f6900000000000000000000000000000000000000000000
cd2000004eab00004c2c00000000000000000000000000000000000000000000
cb380000502400004dc700000000000000000000000000000000000000000000
c843000050c900004f2900000000000000000000000000000000000000000000
d0f8000048ae0000388100000000000000000000000000000000000000000000
d01c00004c2b000047d900000000000000000000000000000000000000000000
ce7200004df000004b7800000000000000000000000000000000000000000000
d31d0000c4ab0000ca9f00000000000000000000000000000000000000000000
d2ef0000c1900000c9b000000000000000000000000000000000000000000000
d2990000ae9a0000c85900000000000000000000000000000000000000000000
d3c90000c46c0000cafd00000000000000000000000000000000000000000000
d40f0000c57f0000cb8a00000000000000000000000000000000000000000000
d4050000c5660000caf000000000000000000000000000000000000000000000
d318000045c30000c43900000000000000000000000000000000000000000000
d338000046240000c3bd00000000000000000000000000000000000000000000
d373000044f20000c35700000000000000000000000000000000000000000000
d29d0000497800003dfb00000000000000000000000000000000000000000000
d24d00004af60000447400000000000000000000000000000000000000000000
d2f8000048370000ac4a00000000000000000000000000000000000000000000
d27800004c56000047d300000000000000000000000000000000000000000000
d1ad00004dcc00004ad400000000000000000000000000000000000000000000
d29400004b440000457200000000000000000000000000000000000000000000
d3b600004e1b00004a3200000000000000000000000000000000000000000000
d28100004fd000004ceb00000000000000000000000000000000000000000000
d32100004dad000049d100000000000000000000000000000000000000000000
d4ac00004db80000487600000000000000000000000000000000000000000000
d43b00004ece00004ad900000000000000000000000000000000000000000000
d42100004dbe0000493600000000000000000000000000000000000000000000
d47d00004bc50000421800000000000000000000000000000000000000000000
d4b6000049170000bf8200000000000000000000000000000000000000000000
d472000049040000be1300000000000000000000000000000000000000000000
d3370000497b00003da100000000000000000000000000000000000000000000
d4a40000c8000000cc2600000000000000000000000000000000000000000000
d48a0000c7e60000cc1e00000000000000000000000000000000000000000000
cf9800004d8600004bbe00000000000000000000000000000000000000000000
d3220000c45b0000c97300000000000000000000000000000000000000000000
d4290000caf30000cd1c00000000000000000000000000000000000000000000
c8250000504a00004f5400000000000000000000000000000000000000000000
cdc500004d9900004c3600000000000000000000000000000000000000000000
d13c0000441b0000bdd000000000000000000000000000000000000000000000
c94900004fee00004ead00000000000000000000000000000000000000000000
c4be0000510a0000505c00000000000000000000000000000000000000000000
cc3d00004f7d00004dea00000000000000000000000000000000000000000000
d02b00004acb0000481300000000000000000000000000000000000000000000
cb2b0000505500004f2b00000000000000000000000000000000000000000000
c9fa0000510000004fe900000000000000000000000000000000000000000000
d3370000c4c40000ca0000000000000000000000000000000000000000000000
d150000049740000435200000000000000000000000000000000000000000000
cdd000004ff700004dba00000000000000000000000000000000000000000000
d3890000bcf60000c95000000000000000000000000000000000000000000000
d42e0000c7bf0000cc4a00000000000000000000000000000000000000000000
d1ca00004a070000414b00000000000000000000000000000000000000000000
d3dd000044610000c65e00000000000000000000000000000000000000000000
d3a1000045690000c4fe00000000000000000000000000000000000000000000
d2e20000478f0000c0ed00000000000000000000000000000000000000000000
d437000044920000c70800000000000000000000000000000000000000000000
d40c000045db0000c52b00000000000000000000000000000000000000000000
d3de00003d050000c86500000000000000000000000000000000000000000000
d47f0000c5690000cc3000000000000000000000000000000000000000000000
d4540000c3ae0000cb1400000000000000000000000000000000000000000000
d3f60000c0060000c9d800000000000000000000000000000000000000000000
d3b10000c4610000cba900000000000000000000000000000000000000000000
d3e60000c63c0000cba400000000000000000000000000000000000000000000
d32f0000b1f00000c84300000000000000000000000000000000000000000000
d30a0000c0320000c93700000000000000000000000000000000000000000000
d3350000c0a30000c92b00000000000000000000000000000000000000000000
d29b000042480000c32a00000000000000000000000000000000000000000000
d2b9000042a60000c17500000000000000000000000000000000000000000000
d2a6000045ba0000357f00000000000000000000000000000000000000000000
d1eb000049cd0000463b00000000000000000000000000000000000000000000
d28100004a200000481d00000000000000000000000000000000000000000000
d1b800004ce900004bd200000000000000000000000000000000000000000000
d0f600004e6e00004d6d00000000000000000000000000000000000000000000
d34800004aa3000048eb00000000000000000000000000000000000000000000
d1b900004eec00004e1100000000000000000000000000000000000000000000
d0d3000050700000500200000000000000000000000000000000000000000000
d2c600004d7600004d2900000000000000000000000000000000000000000000
d148000050550000501e00000000000000000000000000000000000000000000
d1300000507f0000505000000000000000000000000000000000000000000000
d2b600004dc400004e0100000000000000000000000000000000000000000000
d10d000050a40000509600000000000000000000000000000000000000000000
d055000051180000511700000000000000000000000000000000000000000000
d1d500004f6600004fa300000000000000000000000000000000000000000000
d087000050e50000510400000000000000000000000000000000000000000000
d00c0000514f0000515000000000000000000000000000000000000000000000
d1a000004f7100004f9e00000000000000000000000000000000000000000000
d091000050cb000050e300000000000000000000000000000000000000000000
d0020000511b0000511c00000000000000000000000000000000000000000000
d0da000050770000506700000000000000000000000000000000000000000000
cf2a0000519e0000518f00000000000000000000000000000000000000000000
d09a000050530000504b00000000000000000000000000000000000000000000
d16d00004f6000004eb500000000000000000000000000000000000000000000
cfe10000513f000050ea00000000000000000000000000000000000000000000
d037000050a90000506d00000000000000000000000000000000000000000000
d19300004df300004c9800000000000000000000000000000000000000000000
d0c400004fb300004e5900000000000000000000000000000000000000000000
d0640000502200004ee900000000000000000000000000000000000000000000
d1e400004baa000047c400000000000000000000000000000000000000000000
d16300004cec00004a3f00000000000000000000000000000000000000000000
d14300004d2b00004abd00000000000000000000000000000000000000000000
d05b00004e8000004c0100000000000000000000000000000000000000000000
cf190000500400004df000000000000000000000000000000000000000000000
d0ab00004de000004b9200000000000000000000000000000000000000000000
cd330000510700004fa300000000000000000000000000000000000000000000
cd3d0000511b00004fc100000000000000000000000000000000000000000000
d09300004eca00004c5400000000000000000000000000000000000000000000
cad60000520a0000513000000000000000000000000000000000000000000000
ce95000050c400004f9d00000000000000000000000000000000000000000000
d12600004e6200004c6d00000000000000000000000000000000000000000000
ce62000050b7000050c200000000000000000000000000000000000000000000
cf8b000050710000507900000000000000000000000000000000000000000000
d034000050840000506900000000000000000000000000000000000000000000
ce43000051200000517a00000000000000000000000000000000000000000000
cfd1000050a9000050e900000000000000000000000000000000000000000000
cfcb000051480000514a00000000000000000000000000000000000000000000
cd7f000051c80000520600000000000000000000000000000000000000000000
ceac0000517b000051ba00000000000000000000000000000000000000000000
ce44000052440000524500000000000000000000000000000000000000000000
ce50000051e00000521b00000000000000000000000000000000000000000000
ce2e000052030000523f00000000000000000000000000000000000000000000
ce23000052570000525900000000000000000000000000000000000000000000
cdcd000052b2000052d000000000000000000000000000000000000000000000
cd7c000052e80000530700000000000000000000000000000000000000000000
ccc8000053040000530400000000000000000000000000000000000000000000
cf63000051e20000520000000000000000000000000000000000000000000000
cd46000052be000052e000000000000000000000000000000000000000000000
c86a000054010000540200000000000000000000000000000000000000000000
cc30000053440000536200000000000000000000000000000000000000000000
cd100000524b0000528700000000000000000000000000000000000000000000
cb52000052570000527900000000000000000000000000000000000000000000
cd1f000053120000532c00000000000000000000000000000000000000000000
ce9b000051e8000051e700000000000000000000000000000000000000000000
cdae000051070000514400000000000000000000000000000000000000000000
d131000051450000510400000000000000000000000000000000000000000000
d0e400005109000050e700000000000000000000000000000000000000000000
d07b0000501c0000503800000000000000000000000000000000000000000000
d1a5000050cb0000508a00000000000000000000000000000000000000000000
d13e0000508c0000504c00000000000000000000000000000000000000000000
ce9d000051420000512200000000000000000000000000000000000000000000
cf60000051290000510700000000000000000000000000000000000000000000
d01e0000506f0000504e00000000000000000000000000000000000000000000
cd5a000050c7000050e400000000000000000000000000000000000000000000
cf600000508c0000502c00000000000000000000000000000000000000000000
cfbf0000502e00004f9c00000000000000000000000000000000000000000000
ce4a0000502c00004fd800000000000000000000000000000000000000000000
cf9e00004f6200004ede00000000000000000000000000000000000000000000
cffc00004f5d00004e6000000000000000000000000000000000000000000000
cff600004f5b00004e5e00000000000000000000000000000000000000000000
cb1f00005139000050da00000000000000000000000000000000000000000000
cebb0000500e00004ea300000000000000000000000000000000000000000000
d05400004f2000004d6800000000000000000000000000000000000000000000
cc1c000050b20000501500000000000000000000000000000000000000000000
cfdc00004ef300004d7400000000000000000000000000000000000000000000
d1a000004d7800004b7400000000000000000000000000000000000000000000
cbd4000051210000506300000000000000000000000000000000000000000000
cec50000504100004f0200000000000000000000000000000000000000000000
d20300004de400004aef00000000000000000000000000000000000000000000
cf1c0000509600004efc00000000000000000000000000000000000000000000
d14d00004f0400004c9800000000000000000000000000000000000000000000
d2e100004d6d0000496700000000000000000000000000000000000000000000
d1d600004dea00004ae200000000000000000000000000000000000000000000
d32e00004b66000044c900000000000000000000000000000000000000000000
d42a000049470000b6c900000000000000000000000000000000000000000000
d3b8000048860000bb7d00000000000000000000000000000000000000000000
d4130000463c0000c38e00000000000000000000000000000000000000000000
d43f000044060000c61600000000000000000000000000000000000000000000
d2d000004c120000464c00000000000000000000000000000000000000000000
d26200004c6c0000484500000000000000000000000000000000000000000000
d30b0000495200003e0c00000000000000000000000000000000000000000000
d1ce00004d020000497500000000000000000000000000000000000000000000
d0f200004e5500004c1400000000000000000000000000000000000000000000
d18d00004c360000485600000000000000000000000000000000000000000000
d1fe00004c0a0000472c00000000000000000000000000000000000000000000
d1b800004c3a0000485f00000000000000000000000000000000000000000000
d2020000481a00003c1200000000000000000000000000000000000000000000
d4200000c5800000cad300000000000000000000000000000000000000000000
d3c80000c4160000c9a300000000000000000000000000000000000000000000
d3820000c7e10000cb0a00000000000000000000000000000000000000000000
d41f0000c91b0000cc5800000000000000000000000000000000000000000000
d3840000c6140000ca8c00000000000000000000000000000000000000000000
d3570000c8740000cb7a00000000000000000000000000000000000000000000
d3590000c6510000c9d900000000000000000000000000000000000000000000
d37a0000c8090000cab900000000000000000000000000000000000000000000
d4060000cab20000ccd800000000000000000000000000000000000000000000
d2aa0000c06e0000c73b00000000000000000000000000000000000000000000
d3ae0000c8a80000cb2900000000000000000000000000000000000000000000
d4680000cc670000ce1700000000000000000000000000000000000000000000
d177000047350000448c00000000000000000000000000000000000000000000
d2bc0000c0af0000c4fb00000000000000000000000000000000000000000000
d45e0000cac60000ccea00000000000000000000000000000000000000000000
d0b200004bd600004a6e00000000000000000000000000000000000000000000
d19b0000492c0000478e00000000000000000000000000000000000000000000
d36d00003af30000c50900000000000000000000000000000000000000000000
d01500004e7300004de100000000000000000000000000000000000000000000
d09a00004dd600004d4600000000000000000000000000000000000000000000
d19100004cc000004b4c00000000000000000000000000000000000000000000
d00800004fa700004ef500000000000000000000000000000000000000000000
d05e00004f8700004ed700000000000000000000000000000000000000000000
d0a600004fb400004e8800000000000000000000000000000000000000000000
d0b400004f4900004e8800000000000000000000000000000000000000000000
d0d500004f4900004e8800000000000000000000000000000000000000000000
d10c00004f6800004e2c00000000000000000000000000000000000000000000
d17800004ebb00004dcb00000000000000000000000000000000000000000000
d11900004f4200004e5300000000000000000000000000000000000000000000
d18200004e9000004d5200000000000000000000000000000000000000000000
d10e00004fd500004ed300000000000000000000000000000000000000000000
d0c60000503200004f6400000000000000000000000000000000000000000000
d0910000503c00004f3800000000000000000000000000000000000000000000
d1110000508300004fd900000000000000000000000000000000000000000000
d0e40000509800004fd600000000000000000000000000000000000000000000
d0a80000509400004fbc00000000000000000000000000000000000000000000
d25e0000506800004ee200000000000000000000000000000000000000000000
d2490000505400004ecf00000000000000000000000000000000000000000000
d1d50000501f00004e9000000000000000000000000000000000000000000000
d2eb0000504a00004e5600000000000000000000000000000000000000000000
d2770000506b00004ed400000000000000000000000000000000000000000000
d2180000501800004e6e00000000000000000000000000000000000000000000
d2190000500c00004e5600000000000000000000000000000000000000000000
d1c30000504b00004ee900000000000000000000000000000000000000000000
d19800004fdd00004e4600000000000000000000000000000000000000000000
d0f400004fad00004e5600000000000000000000000000000000000000000000
d08a0000505200004f4d00000000000000000000000000000000000000000000
d0a500004f9e00004e6f00000000000000000000000000000000000000000000
cfb300004f6e00004e0500000000000000000000000000000000000000000000
cc9600005156000050a100000000000000000000000000000000000000000000
caf6000051ad0000513f00000000000000000000000000000000000000000000
cc1d000050ab00004ffd00000000000000000000000000000000000000000000
c1b00000526d000051c000000000000000000000000000000000000000000000
41860000533b000052d800000000000000000000000000000000000000000000
c9b8000051360000509500000000000000000000000000000000000000000000
40aa000052fc0000525c00000000000000000000000000000000000000000000
470d000053d10000536f00000000000000000000000000000000000000000000
cd11000050b80000500500000000000000000000000000000000000000000000
c75400005265000051b200000000000000000000000000000000000000000000
beb0000053330000529900000000000000000000000000000000000000000000
d06a00004f1b00004d2b00000000000000000000000000000000000000000000
cdbc000051170000504400000000000000000000000000000000000000000000
cb9b0000520e0000513b00000000000000000000000000000000000000000000
d12900004ed500004c7200000000000000000000000000000000000000000000
cee5000051250000500e00000000000000000000000000000000000000000000
cc61000052560000516200000000000000000000000000000000000000000000
d03b000050b000004ee100000000000000000000000000000000000000000000
ce44000051da0000509a00000000000000000000000000000000000000000000
cc80000052ae0000518a00000000000000000000000000000000000000000000
ce75000051be0000507f00000000000000000000000000000000000000000000
ce24000051f9000050b900000000000000000000000000000000000000000000
cdf400005232000050f200000000000000000000000000000000000000000000
cf740000512e00004fdd00000000000000000000000000000000000000000000
cf0c000051840000504400000000000000000000000000000000000000000000
cee3000051e70000508600000000000000000000000000000000000000000000
d0c00000504a00004e1400000000000000000000000000000000000000000000
d0450000511700004f8d00000000000000000000000000000000000000000000
d0350000518400004fec00000000000000000000000000000000000000000000
d15d0000506a00004e1600000000000000000000000000000000000000000000
d0e20000510800004f4f00000000000000000000000000000000000000000000
d11e000050dc00004eba00000000000000000000000000000000000000000000
d1ad000050c900004e9300000000000000000000000000000000000000000000
d151000050fb00004f1500000000000000000000000000000000000000000000
d123000050cb00004ed300000000000000000000000000000000000000000000
d18f0000508000004e5c00000000000000000000000000000000000000000000
d19e0000506300004e2100000000000000000000000000000000000000000000
d104000050bc00004ef200000000000000000000000000000000000000000000
d0be0000509d00004efb00000000000000000000000000000000000000000000
d0e20000508b00004ed600000000000000000000000000000000000000000000
d0ac000050c100004f4200000000000000000000000000000000000000000000
cf18000051ac0000508d00000000000000000000000000000000000000000000
cf30000051b30000509200000000000000000000000000000000000000000000
d02a000051210000500100000000000000000000000000000000000000000000
ce070000520c000050fa00000000000000000000000000000000000000000000
ce7d000051e2000050d000000000000000000000000000000000000000000000
cf99000051550000504200000000000000000000000000000000000000000000
ce18000051c0000050c000000000000000000000000000000000000000000000
ceb20000515d0000506900000000000000000000000000000000000000000000
cdb2000051b5000050a800000000000000000000000000000000000000000000
cca9000052240000513100000000000000000000000000000000000000000000
cd0e000051a4000050b700000000000000000000000000000000000000000000
c97f0000523b0000513500000000000000000000000000000000000000000000
c6af000052e00000520000000000000000000000000000000000000000000000
c313000052ea000051f700000000000000000000000000000000000000000000
465c0000530f0000524700000000000000000000000000000000000000000000
2f1b000053070000522700000000000000000000000000000000000000000000
44e90000531a0000524600000000000000000000000000000000000000000000
4de6000053e20000534000000000000000000000000000000000000000000000
46a0000053b0000052d000000000000000000000000000000000000000000000
48530000532c0000526b00000000000000000000000000000000000000000000
50f7000054a10000545000000000000000000000000000000000000000000000
4828000053fd0000531d00000000000000000000000000000000000000000000
4a0c0000538a000052c900000000000000000000000000000000000000000000
525c00005532000054ec00000000000000000000000000000000000000000000
48450000541c0000538300000000000000000000000000000000000000000000
48300000535c000052a700000000000000000000000000000000000000000000
52b70000557f0000554900000000000000000000000000000000000000000000
45eb000053f90000539800000000000000000000000000000000000000000000
4974000053e10000536100000000000000000000000000000000000000000000
51bb000055400000550400000000000000000000000000000000000000000000
481900005412000053eb00000000000000000000000000000000000000000000
4a18000053e1000053b400000000000000000000000000000000000000000000
502b000054aa0000547b00000000000000000000000000000000000000000000
473c000053ea0000540400000000000000000000000000000000000000000000
4b22000054180000541d00000000000000000000000000000000000000000000
4bf60000538a0000533600000000000000000000000000000000000000000000
c400000053530000537a00000000000000000000000000000000000000000000
4599000054080000541800000000000000000000000000000000000000000000
46ef000053560000533400000000000000000000000000000000000000000000
cc9c000052e00000531500000000000000000000000000000000000000000000
cabc000052f40000530b00000000000000000000000000000000000000000000
bed7000053710000538800000000000000000000000000000000000000000000
cebd000052400000525600000000000000000000000000000000000000000000
ccf1000052b5000052b500000000000000000000000000000000000000000000
c9ab000052c8000052c800000000000000000000000000000000000000000000
cdc3000052570000524e00000000000000000000000000000000000000000000
cdb1000052340000522b00000000000000000000000000000000000000000000
cae8000052700000525900000000000000000000000000000000000000000000
cd5100005204000051ea00000000000000000000000000000000000000000000
c8e10000534e0000531f00000000000000000000000000000000000000000000
c87b000052d30000527b00000000000000000000000000000000000000000000
c8c3000052cd000052be00000000000000000000000000000000000000000000
c6100000533b000052d500000000000000000000000000000000000000000000
3e7d000053b50000536c00000000000000000000000000000000000000000000
c6e9000052d20000528400000000000000000000000000000000000000000000
3c38000053ec0000536d00000000000000000000000000000000000000000000
43b6000053de0000537600000000000000000000000000000000000000000000
c921000052c50000523e00000000000000000000000000000000000000000000
3336000053f20000536000000000000000000000000000000000000000000000
ba02000053ad0000531a00000000000000000000000000000000000000000000
c7360000538a000052d800000000000000000000000000000000000000000000
c7cf00005388000052a300000000000000000000000000000000000000000000
c58c0000539e000052b800000000000000000000000000000000000000000000
ccd00000526c0000516c00000000000000000000000000000000000000000000
cc2e000052d4000051d300000000000000000000000000000000000000000000
ca93000053560000524b00000000000000000000000000000000000000000000
ccbe0000523c0000513700000000000000000000000000000000000000000000
cc9c000052830000517e00000000000000000000000000000000000000000000
cc6400005301000051cd00000000000000000000000000000000000000000000
38ab000053ed000052d700000000000000000000000000000000000000000000
c7ae000053380000521d00000000000000000000000000000000000000000000
c9ef0000532b0000522e00000000000000000000000000000000000000000000
44390000538a000052b300000000000000000000000000000000000000000000
4644000054180000533d00000000000000000000000000000000000000000000
46c200005451000053d200000000000000000000000000000000000000000000
4bc80000542a000053b200000000000000000000000000000000000000000000
4b5700005434000053c700000000000000000000000000000000000000000000
4a360000544a0000541900000000000000000000000000000000000000000000
41bc000052f00000524c00000000000000000000000000000000000000000000
491a000054100000537d00000000000000000000000000000000000000000000
4a38000054540000542100000000000000000000000000000000000000000000
c184000053150000525100000000000000000000000000000000000000000000
c618000052b6000051fc00000000000000000000000000000000000000000000
c94900005257000051da00000000000000000000000000000000000000000000
cdf1000051240000504e00000000000000000000000000000000000000000000
ceff000050910000501100000000000000000000000000000000000000000000
cef70000503a00004fea00000000000000000000000000000000000000000000
ce6d00005104000050a300000000000000000000000000000000000000000000
cf14000050bd0000505d00000000000000000000000000000000000000000000
ce7a000050ca0000506c00000000000000000000000000000000000000000000
caee000052770000521a00000000000000000000000000000000000000000000
ccb3000051ae0000515200000000000000000000000000000000000000000000
cd95000050e2000050a000000000000000000000000000000000000000000000
cca5000051440000514400000000000000000000000000000000000000000000
cc42000051850000518600000000000000000000000000000000000000000000
ca2400005200000051c200000000000000000000000000000000000000000000
cca2000050ca000050e800000000000000000000000000000000000000000000
cc3a0000510c0000512c00000000000000000000000000000000000000000000
cb770000516a0000512f00000000000000000000000000000000000000000000
cc20000050cb000050ea00000000000000000000000000000000000000000000
c9f90000516c0000518c00000000000000000000000000000000000000000000
c87a000051cb000051eb00000000000000000000000000000000000000000000
c85400005168000051a600000000000000000000000000000000000000000000
3a4a000052a4000052e400000000000000000000000000000000000000000000
44d5000053260000536500000000000000000000000000000000000000000000
c6af000051a70000520400000000000000000000000000000000000000000000
44b7000053220000538100000000000000000000000000000000000000000000
4866000053a4000053e500000000000000000000000000000000000000000000
c84b000051a80000520600000000000000000000000000000000000000000000
44bd00005361000053c000000000000000000000000000000000000000000000
48e6000054100000542200000000000000000000000000000000000000000000
c3c40000527d000052db00000000000000000000000000000000000000000000
c58000005258000052b800000000000000000000000000000000000000000000
c5580000525e000052bc00000000000000000000000000000000000000000000
cc700000513c0000517c00000000000000000000000000000000000000000000
cb4800005194000051d600000000000000000000000000000000000000000000
cbb600005178000051b900000000000000000000000000000000000000000000
ce7f000050950000509800000000000000000000000000000000000000000000
cddc000050f4000050f800000000000000000000000000000000000000000000
ce8a000050630000506700000000000000000000000000000000000000000000
cdb8000051390000513800000000000000000000000000000000000000000000
ceab000050960000509600000000000000000000000000000000000000000000
cf6a00004fef00004fef00000000000000000000000000000000000000000000
cb3a000052120000521100000000000000000000000000000000000000000000
ceb0000050930000509300000000000000000000000000000000000000000000
ced2000050440000504400000000000000000000000000000000000000000000
cc11000051d2000051d100000000000000000000000000000000000000000000
ceea000050760000507500000000000000000000000000000000000000000000
ce1d0000509f0000509e00000000000000000000000000000000000000000000
cdad000050cc000050cb00000000000000000000000000000000000000000000
ce8b0000506d0000506d00000000000000000000000000000000000000000000
cea8000050570000505700000000000000000000000000000000000000000000
cef60000502000004fcf00000000000000000000000000000000000000000000
ce4c000050850000508300000000000000000000000000000000000000000000
cf9300004fc300004fc200000000000000000000000000000000000000000000
cddb000050ad0000506c00000000000000000000000000000000000000000000
cf7f00004fd700004f6900000000000000000000000000000000000000000000
cf550000500000004f9300000000000000000000000000000000000000000000
ce790000507a0000500300000000000000000000000000000000000000000000
ce7d000050870000501100000000000000000000000000000000000000000000
ced2000050430000500100000000000000000000000000000000000000000000
cf7300004fce00004f3500000000000000000000000000000000000000000000
cd77000050f5000050aa00000000000000000000000000000000000000000000
ce1c0000506a0000507600000000000000000000000000000000000000000000
cf3800004ffe00004f7c00000000000000000000000000000000000000000000
cc180000519f0000515f00000000000000000000000000000000000000000000
cc2b000051570000517400000000000000000000000000000000000000000000
cfec00004f1800004e9500000000000000000000000000000000000000000000
ccd000005129000050e900000000000000000000000000000000000000000000
c9a3000051d2000051ee00000000000000000000000000000000000000000000
d07300004dac00004d2a00000000000000000000000000000000000000000000
cf0100004fb000004f2f00000000000000000000000000000000000000000000
cc5c000050fe0000511b00000000000000000000000000000000000000000000
ce9e00004f4600004f5700000000000000000000000000000000000000000000
ce5800004fa900004fbd00000000000000000000000000000000000000000000
ccfe00005063000050b200000000000000000000000000000000000000000000
cc300000507c000050b200000000000000000000000000000000000000000000
cc490000507d000050b500000000000000000000000000000000000000000000
cb04000050d90000513800000000000000000000000000000000000000000000
c9d1000050d90000511700000000000000000000000000000000000000000000
c945000051390000517800000000000000000000000000000000000000000000
c4040000520a0000526900000000000000000000000000000000000000000000
cb800000508c000050ca00000000000000000000000000000000000000000000
c947000051390000517800000000000000000000000000000000000000000000
c00f00005277000052d600000000000000000000000000000000000000000000
ccdd0000500f0000504d00000000000000000000000000000000000000000000
caa4000051260000514f00000000000000000000000000000000000000000000
c38a00005252000052b000000000000000000000000000000000000000000000
cd7e0000502f0000505600000000000000000000000000000000000000000000
ccc0000050b7000050d700000000000000000000000000000000000000000000
cb090000514d0000517e00000000000000000000000000000000000000000000
cfb400004f3400004eec00000000000000000000000000000000000000000000
cf00000050040000500c00000000000000000000000000000000000000000000
ce18000050780000508100000000000000000000000000000000000000000000
cf6f0000505000004ff200000000000000000000000000000000000000000000
cf940000504e0000500c00000000000000000000000000000000000000000000
cf46000050360000503300000000000000000000000000000000000000000000
cf0b000051090000509300000000000000000000000000000000000000000000
cf54000050cd0000506c00000000000000000000000000000000000000000000
cf7f000050590000505600000000000000000000000000000000000000000000
ce51000051910000511000000000000000000000000000000000000000000000
ce6e00005155000050f400000000000000000000000000000000000000000000
ce5c00005100000050fc00000000000000000000000000000000000000000000
ccc5000051f1000051c100000000000000000000000000000000000000000000
cd300000518d0000516a00000000000000000000000000000000000000000000
cc57000051b0000051ae00000000000000000000000000000000000000000000
cd65000051180000511600000000000000000000000000000000000000000000
cd61000050eb000050ff00000000000000000000000000000000000000000000
cb6e000051a8000051bc00000000000000000000000000000000000000000000
cc75000050ec000050fe00000000000000000000000000000000000000000000
ccab000050c7000050e600000000000000000000000000000000000000000000
cb440000514b0000516b00000000000000000000000000000000000000000000
cbb3000050b6000050e800000000000000000000000000000000000000000000
c7bb000051ba000051ed00000000000000000000000000000000000000000000
be560000527e000052b100000000000000000000000000000000000000000000
c87f0000515d0000519b00000000000000000000000000000000000000000000
455c000053360000537600000000000000000000000000000000000000000000
4a9a000054060000542600000000000000000000000000000000000000000000
4013000052f50000532100000000000000000000000000000000000000000000
496a0000540e0000542500000000000000000000000000000000000000000000
4aa80000540e0000542e00000000000000000000000000000000000000000000
4407000053c8000053d500000000000000000000000000000000000000000000
4677000054010000541100000000000000000000000000000000000000000000
42b8000053530000538000000000000000000000000000000000000000000000
c785000052f0000052ef00000000000000000000000000000000000000000000
c5ce000052f90000530600000000000000000000000000000000000000000000
c883000052520000526000000000000000000000000000000000000000000000
ccb2000051c1000051c000000000000000000000000000000000000000000000
ccfc000051900000519000000000000000000000000000000000000000000000
cd16000051650000516500000000000000000000000000000000000000000000
ce6d000050e4000050e200000000000000000000000000000000000000000000
cf23000050990000509900000000000000000000000000000000000000000000
cea9000050d6000050d600000000000000000000000000000000000000000000
cf600000502a0000500800000000000000000000000000000000000000000000
cf5e0000503b0000501a00000000000000000000000000000000000000000000
cf04000050870000508600000000000000000000000000000000000000000000
cec30000500b00004f9300000000000000000000000000000000000000000000
cec00000503a00004ff400000000000000000000000000000000000000000000
cee00000505a0000505700000000000000000000000000000000000000000000
cd4c000050490000501800000000000000000000000000000000000000000000
ce1f0000502d00004ff800000000000000000000000000000000000000000000
ced90000502c0000500c00000000000000000000000000000000000000000000
caed000050c4000050a200000000000000000000000000000000000000000000
cd030000504a0000502900000000000000000000000000000000000000000000
ce7c000050470000500700000000000000000000000000000000000000000000
c37e000051e5000051b600000000000000000000000000000000000000000000
ca5b00005121000050e400000000000000000000000000000000000000000000
cceb000050f2000050b200000000000000000000000000000000000000000000
47ad00005361000052f600000000000000000000000000000000000000000000
c4a500005235000051b800000000000000000000000000000000000000000000
ca44000051b60000516600000000000000000000000000000000000000000000
498a000053ed0000533100000000000000000000000000000000000000000000
3816000052e80000522c00000000000000000000000000000000000000000000
c6580000526f000051e400000000000000000000000000000000000000000000
4698000053630000527500000000000000000000000000000000000000000000
3d21000053050000520b00000000000000000000000000000000000000000000
c16a000052d20000520200000000000000000000000000000000000000000000
4857000053530000526c00000000000000000000000000000000000000000000
4379000053010000520700000000000000000000000000000000000000000000
b918000052d30000520b00000000000000000000000000000000000000000000
4a3f000053b8000052eb00000000000000000000000000000000000000000000
46c9000053290000527400000000000000000000000000000000000000000000
ac38000052c30000521600000000000000000000000000000000000000000000
3a1b000053390000527d00000000000000000000000000000000000000000000
c5290000529a000051f900000000000000000000000000000000000000000000
caef000051e40000513100000000000000000000000000000000000000000000
cc4200005270000051d800000000000000000000000000000000000000000000
cdcf000051e00000513400000000000000000000000000000000000000000000
cf45000051250000507900000000000000000000000000000000000000000000
cf540000520f0000515a00000000000000000000000000000000000000000000
d04200005162000050ad00000000000000000000000000000000000000000000
d0960000510d0000505800000000000000000000000000000000000000000000
d04f000051a80000510800000000000000000000000000000000000000000000
d107000051040000506400000000000000000000000000000000000000000000
d10b000051000000505f00000000000000000000000000000000000000000000
cec500005219000051a200000000000000000000000000000000000000000000
d07500005124000050ad00000000000000000000000000000000000000000000
d0a30000510a0000509300000000000000000000000000000000000000000000
c95900005306000052ee00000000000000000000000000000000000000000000
cd30000051eb000051d400000000000000000000000000000000000000000000
cdfc000051cd000051ad00000000000000000000000000000000000000000000
c852000053060000530400000000000000000000000000000000000000000000
c987000052e5000052db00000000000000000000000000000000000000000000
c9e600005318000052f900000000000000000000000000000000000000000000
c973000052f4000052e900000000000000000000000000000000000000000000
c913000053600000534000000000000000000000000000000000000000000000
c9360000536f0000534f00000000000000000000000000000000000000000000
ccd2000052ac0000528200000000000000000000000000000000000000000000
cbc1000053370000530e00000000000000000000000000000000000000000000
cb8d000053330000530a00000000000000000000000000000000000000000000
cea1000052670000522600000000000000000000000000000000000000000000
cda6000052f8000052b800000000000000000000000000000000000000000000
cc8a00005338000052f800000000000000000000000000000000000000000000
cdf6000052860000524d00000000000000000000000000000000000000000000
cdb3000052ab0000527300000000000000000000000000000000000000000000
cc8b000052c30000529200000000000000000000000000000000000000000000
cae10000530b000052e900000000000000000000000000000000000000000000
ccd6000052390000521900000000000000000000000000000000000000000000
ccbd000051c2000051c100000000000000000000000000000000000000000000
c7dd0000537e0000536b00000000000000000000000000000000000000000000
cccf0000521c0000520a00000000000000000000000000000000000000000000
cd7b0000514d0000515300000000000000000000000000000000000000000000
c7a0000053720000539000000000000000000000000000000000000000000000
cabc000052af000052cf00000000000000000000000000000000000000000000
cd3c000051ad000051d300000000000000000000000000000000000000000000
c1d30000538c000053ab00000000000000000000000000000000000000000000
c958000052a4000052c300000000000000000000000000000000000000000000
cc07000051a0000051d800000000000000000000000000000000000000000000
3f94000053310000535500000000000000000000000000000000000000000000
c4160000527a000052a000000000000000000000000000000000000000000000
c74c000051e10000520600000000000000000000000000000000000000000000
49b00000538f000053c300000000000000000000000000000000000000000000
45c6000052cf0000530400000000000000000000000000000000000000000000
3fbf0000523a0000528400000000000000000000000000000000000000000000
4da7000054390000543800000000000000000000000000000000000000000000
4bd6000053920000539600000000000000000000000000000000000000000000
4a9a000052b10000531f00000000000000000000000000000000000000000000
4df0000054590000545300000000000000000000000000000000000000000000
4de60000542b0000543800000000000000000000000000000000000000000000
4e67000054180000542700000000000000000000000000000000000000000000
4a3a0000540a000053cb00000000000000000000000000000000000000000000
4cb0000054350000542e00000000000000000000000000000000000000000000
4efb000054750000548200000000000000000000000000000000000000000000
c9000000527b000051f700000000000000000000000000000000000000000000
35090000533f000052d700000000000000000000000000000000000000000000
49f3000053d6000053cc00000000000000000000000000000000000000000000
d0b80000502100004ef500000000000000000000000000000000000000000000
ceff000051030000506600000000000000000000000000000000000000000000
cc700000516a0000512d00000000000000000000000000000000000000000000
d21100004fde00004e2300000000000000000000000000000000000000000000
d0500000510c0000508700000000000000000000000000000000000000000000
cd42000051a40000519d00000000000000000000000000000000000000000000
d0d50000517b000050bd00000000000000000000000000000000000000000000
ce79000052ae0000521400000000000000000000000000000000000000000000
cc10000052eb000052c700000000000000000000000000000000000000000000
ceec00005276000051db00000000000000000000000000000000000000000000
cd270000532b000052eb00000000000000000000000000000000000000000000
cb820000530a000052ec00000000000000000000000000000000000000000000
cb2a000053610000532300000000000000000000000000000000000000000000
c9fa000053650000534700000000000000000000000000000000000000000000
c9f5000052ea0000530b00000000000000000000000000000000000000000000
c83d000053000000530100000000000000000000000000000000000000000000
c8d6000052ea0000530b00000000000000000000000000000000000000000000
c8e30000528f000052ed00000000000000000000000000000000000000000000
c33b00005246000052a400000000000000000000000000000000000000000000
bbbe000052ab0000530a00000000000000000000000000000000000000000000
c1b9000052ab0000532a00000000000000000000000000000000000000000000
bd82000051e50000526000000000000000000000000000000000000000000000
4074000052c20000532100000000000000000000000000000000000000000000
35d6000052a70000534300000000000000000000000000000000000000000000
*/

	end
`endif
`ifdef SACC
	reg [169*16-1:0] avepooldata;
	initial begin
		avepooldata = {16'h3757, 16'h39da, 16'h3b67, 16'h3376, 16'h3bb5, 16'h30da, 16'h3b8a, 16'h2675, 16'h3454, 16'h2d3e, 16'h39d1, 16'h3614, 16'h36dd,
	16'h304e, 16'h3023, 16'h3b02, 16'h3367, 16'h3b9d, 16'h32ff, 16'h387e, 16'h384d, 16'h3812, 16'h3bad, 16'h3587, 16'h33f5, 16'h3ab1,
	16'h3945, 16'h3625, 16'h2f8f, 16'h39de, 16'h367c, 16'h287c, 16'h354f, 16'h2d21, 16'h39a8, 16'h382e, 16'h3b5c, 16'h3ba0, 16'h39cd,
	16'h3a0c, 16'h2e91, 16'h38cb, 16'h2bc9, 16'h3872, 16'h3173, 16'h37b0, 16'h32da, 16'h3b5a, 16'h380e, 16'h3892, 16'h3988, 16'h390d,
	16'h38e9, 16'h3a7c, 16'h3a78, 16'h3a50, 16'h3894, 16'h397d, 16'h314d, 16'h2c73, 16'h304c, 16'h3774, 16'h36ca, 16'h3512, 16'h3b17,
	16'h363f, 16'h3721, 16'h3489, 16'h2fe5, 16'h34c6, 16'h3aaf, 16'h37b1, 16'h38e3, 16'h36e3, 16'h3942, 16'h3bbe, 16'h39ac, 16'h3873,
	16'h37c1, 16'h340b, 16'h3b26, 16'h3b70, 16'h372c, 16'h36f3, 16'h3bd5, 16'h3a3a, 16'h339e, 16'h3821, 16'h33f5, 16'h3858, 16'h3bf0,
	16'h3beb, 16'h3b73, 16'h3a1c, 16'h3a83, 16'h3bb2, 16'h3808, 16'h39c7, 16'h3b72, 16'h39cf, 16'h2a93, 16'h3402, 16'h39d8, 16'h3974,
	16'h3483, 16'h3b46, 16'h3af9, 16'h38ad, 16'h3933, 16'h30de, 16'h305e, 16'h2fdb, 16'h3ad9, 16'h3ad2, 16'h39fa, 16'h2ae8, 16'h32b6,
	16'h3596, 16'h3b5e, 16'h329c, 16'h2da6, 16'h3a5a, 16'h3562, 16'h3a02, 16'h3a38, 16'h354e, 16'h3b19, 16'h3976, 16'h383c, 16'h29d8,
	16'h3a29, 16'h3a08, 16'h3301, 16'h386f, 16'h2a75, 16'h37cf, 16'h3267, 16'h30e1, 16'h3967, 16'h388a, 16'h397b, 16'h3ab4, 16'h3999,
	16'h3899, 16'h378f, 16'h394b, 16'h3554, 16'h3723, 16'h3880, 16'h327a, 16'h3a9b, 16'h383c, 16'h3936, 16'h387d, 16'h34c5, 16'h3782,
	16'h3a3f, 16'h3b8c, 16'h3156, 16'h3ba7, 16'h3b97, 16'h2e65, 16'h3194, 16'h32d6, 16'h3572, 16'h3889, 16'h3aa1, 16'h36d4, 16'h2cc5}; //16'h558f, 16'h3836
	end
`endif
`ifdef SCMP
	reg [9*16-1:0] maxpooldata;
	initial begin
		maxpooldata = {16'h4880, 16'h4400, 16'h4600, 16'h4880, 16'h4200, 16'h4700, 16'h3c00, 16'h4000, 16'h4500}; //9,4,6,8,3,7,1,2,5
	end
`endif

engine engine_(
	.clk					(clk),
//Control signals csb->engine
	.rst					(rst),
	.engine_valid			(engine_valid),
	.op_type				(op_type),
	.stride					(stride),
	.stride2				(stride2),
	.kernel					(kernel),
	.kernel_size			(kernel_size),
	.i_channel				(i_channel),
	.o_channel				(o_channel),
	.i_side					(i_side),
	.o_side					(o_side),
	.bias					(bias),
//Response signals engine->csb
	.gemm_finish			(gemm_finish),
	.engine_ready			(engine_ready),
//Command path engine->dma
	.dma_p0_writes_en		(dma_p0_writes_en),
	.dma_p2_reads_en		(dma_p2_reads_en),
    .dma_p3_reads_en		(dma_p3_reads_en),
//Data path dma->engine
	.dma_p2_ob_data			(dma_p2_ob_data),
	.dma_p3_ob_data			(dma_p3_ob_data),
	.dma_p2_ob_we			(dma_p2_ob_we),
	.dma_p3_ob_we			(dma_p3_ob_we),
	.dma_p0_ib_data			(dma_p0_ib_data)
);

always #5 clk = ~clk;
reg [7:0] count; initial count = 0;
always @(posedge clk) begin
	if(gemm_finish) engine_valid <= 0; // pull down engine_valid after the whole op is done
end

integer m,n,offset;
initial begin
    rst = 1;
    clk = 0;
    m = 0; n = 0; offset = 0;
    engine_valid = 0;
    op_type = 0; stride = 0; stride2 = 0;
	kernel = 0; kernel_size = 0; i_channel = 0; o_channel = 0; i_side = 0; o_side = 0; 
	dma_p2_ob_data = 16'h0000;
	dma_p3_ob_data = 16'h0000;
	dma_p2_ob_we = 0;
	dma_p3_ob_we = 0;
	bias = 16'h0000;
    #20 rst = 1;
    #10 rst = 0;
`ifdef CMAC
    #100 op_type = 1; stride = 2; stride2 = 6;
		//kernel = 3; kernel_size = 9; i_channel = 3; o_channel = 1; i_side = 227; o_side = 113;
		kernel = 3; kernel_size = 9; i_channel = 3; o_channel = 1; i_side = 7; o_side = 4; bias = 16'hA35C;
`endif
`ifdef SCMP
	#100 op_type = 2; stride = 2; stride2 = 6;
		kernel = 3; kernel_size = 9; i_channel = 8; o_channel = 1; i_side = 3; o_side = 1; bias = 16'h0000;
`endif
`ifdef SACC
	#100 op_type = 3; stride = 1; 
		kernel = 13; kernel_size = 169; i_channel = 3; o_channel = 1; i_side = 13; o_side = 1; bias = 16'h0000;
`endif
    #10 engine_valid = 1;
	//#3000 rst = 1;
	//#20 rst = 0;
	//#20 engine_valid = 1;
end

always @(posedge clk) begin
	if(engine_valid) begin
		if(dma_p2_reads_en) begin 
			dma_p2_ob_we <= 1;
`ifdef CMAC
			dma_p2_ob_data <= data[m]; 
			m <= m + 1; 
`endif
`ifdef SCMP
			dma_p2_ob_data <= maxpooldata[m*16 +: 16];
			offset <= offset + 1;
			if(offset == 7) begin
				m <= m + 1;
				offset <= 0;
			end
`endif
`ifdef SACC
			dma_p2_ob_data <= avepooldata[m*16 +: 16];
			offset <= offset + 1;
			if(offset == 7) begin
				m <= m + 1;
				offset <= 0;
			end
`endif
		end else dma_p2_ob_we <= 0;
`ifdef CMAC
		if(dma_p3_reads_en) begin 
			dma_p3_ob_we <= 1;
			dma_p3_ob_data <= weight[n]; 
			n <= n + 1; 
		end else dma_p3_ob_we <= 0;
`endif
	end
end

endmodule