module csb(

);
endmodule