`ifndef __MACROS__
`define __MACROS__
`define BURST_LEN 8
`define CMD_BURST_LEN 3
`define MAX_O_SIDE 128
`define MAX_KERNEL 3
`define MAX_KERNEL_SIZE 9
`endif