module pool (

);

endmodule