module dma(

);

endmodule