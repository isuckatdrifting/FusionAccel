module pool_3x3 (
    input clk,
    input rst_n,
    input im,
    output om,
    input pool_ready,
    output pool_valid
);

endmodule

//TODO: Bitonic Sort Logic for 13x13 pooling