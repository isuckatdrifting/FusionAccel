module top(

);

usb usb_();
endmodule